*
* MAIN CELL: Component pathname : root_element
*
   .MODEL BDC_switch_ideal "label 1"="TE" "control"=1
   .MODEL "Waveguide Crossing" "label 1"="TE" "transmission 1"=0.9954054174 "cross talk 1"=0.0001
   + "transmission 2"=1 "cross talk 2"=0 "reflection 1"=0.001
   + "reflection 2"=0 "label 2"="TM" "orthogonal identifier 1"=1
   + "orthogonal identifier 2"=2
   .MODEL "Straight Waveguide" "excess loss temperature sensitivity 2"=0 "label 1"="TE" "orthogonal identifier 1"=1 
   + "loss 1"=0 "number of taps"=64 "dispersion 1"=0 
   + "effective index temperature sensitivity 2"=0 "effective index 2"=1 length=10u 
   + "group index 2"=1 "orthogonal identifier 2"=2 "nominal temperature"=300 
   + "loss 2"=0 "dispersion 2"=0 frequency=193.1T 
   + "digital filter"=0 "run diagnostic"=0 "window function"="rectangular" 
   + "thermal fill factor"=1 "excess loss temperature sensitivity 1"=0 "label 2"="TM" 
   + "thermal effects"=0 "effective index temperature sensitivity 1"=0 "effective index 1"=1 

.subckt HDBE  N$34561 N$34563 N$34565 N$34567 N$34569 N$34571 N$34573 N$34575 N$34577 N$34579 N$34581 N$34583 N$34585 N$34587 N$34589 N$34591 N$34593 N$34595 N$34597 N$34599 N$34601 N$34603 N$34605 N$34607 N$34609 N$34611 N$34613 N$34615 N$34617 N$34619 N$34621 N$34623 N$34625 N$34627 N$34629 N$34631 N$34633 N$34635 N$34637 N$34639 N$34641 N$34643 N$34645 N$34647 N$34649 N$34651 N$34653 N$34655 N$34657 N$34659 N$34661 N$34663 N$34665 N$34667 N$34669 N$34671 N$34673 N$34675 N$34677 N$34679 N$34681 N$34683 N$34685 N$34687 N$34945 N$34947 N$34949 N$34951 N$34953 N$34955 N$34957 N$34959 N$34961 N$34963 N$34965 N$34967 N$34969 N$34971 N$34973 N$34975 N$34977 N$34979 N$34981 N$34983 N$34985 N$34987 N$34989 N$34991 N$34993 N$34995 N$34997 N$34999 N$35001 N$35003 N$35005 N$35007 N$35009 N$35011 N$35013 N$35015 N$35017 N$35019 N$35021 N$35023 N$35025 N$35027 N$35029 N$35031 N$35033 N$35035 N$35037 N$35039 N$35041 N$35043 N$35045 N$35047 N$35049 N$35051 N$35053 N$35055 N$35057 N$35059 N$35061 N$35063 N$35065 N$35067 N$35069 N$35071
   S4609 N$34561 N$34562 N$26237 N$17922 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4610 N$34563 N$34564 N$17924 N$17926 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4611 N$34565 N$34566 N$17928 N$17930 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4612 N$34567 N$34568 N$17932 N$17934 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4613 N$34569 N$34570 N$17936 N$17938 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4614 N$34571 N$34572 N$17940 N$17942 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4615 N$34573 N$34574 N$17944 N$17946 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4616 N$34575 N$34576 N$17948 N$17950 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4617 N$34577 N$34578 N$17952 N$17954 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4618 N$34579 N$34580 N$17956 N$17958 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4619 N$34581 N$34582 N$17960 N$17962 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4620 N$34583 N$34584 N$17964 N$17966 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4621 N$34585 N$34586 N$17968 N$17970 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4622 N$34587 N$34588 N$17972 N$17974 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4623 N$34589 N$34590 N$17976 N$17978 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4624 N$34591 N$34592 N$17980 N$17982 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4625 N$34593 N$34594 N$17984 N$17986 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4626 N$34595 N$34596 N$17988 N$17990 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4627 N$34597 N$34598 N$17992 N$17994 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4628 N$34599 N$34600 N$17996 N$17998 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4629 N$34601 N$34602 N$18000 N$18002 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4630 N$34603 N$34604 N$18004 N$18006 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4631 N$34605 N$34606 N$18008 N$18010 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4632 N$34607 N$34608 N$18012 N$18014 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4633 N$34609 N$34610 N$18016 N$18018 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4634 N$34611 N$34612 N$18020 N$18022 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4635 N$34613 N$34614 N$18024 N$18026 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4636 N$34615 N$34616 N$18028 N$18030 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4637 N$34617 N$34618 N$18032 N$18034 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4638 N$34619 N$34620 N$18036 N$18038 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4639 N$34621 N$34622 N$18040 N$18042 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4640 N$34623 N$34624 N$18044 N$18046 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4641 N$34625 N$34626 N$18048 N$18050 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4642 N$34627 N$34628 N$18052 N$18054 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4643 N$34629 N$34630 N$18056 N$18058 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4644 N$34631 N$34632 N$18060 N$18062 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4645 N$34633 N$34634 N$18064 N$18066 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4646 N$34635 N$34636 N$18068 N$18070 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4647 N$34637 N$34638 N$18072 N$18074 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4648 N$34639 N$34640 N$18076 N$18078 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4649 N$34641 N$34642 N$18080 N$18082 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4650 N$34643 N$34644 N$18084 N$18086 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4651 N$34645 N$34646 N$18088 N$18090 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4652 N$34647 N$34648 N$18092 N$18094 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4653 N$34649 N$34650 N$18096 N$18098 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4654 N$34651 N$34652 N$18100 N$18102 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4655 N$34653 N$34654 N$18104 N$18106 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4656 N$34655 N$34656 N$18108 N$18110 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4657 N$34657 N$34658 N$18112 N$18114 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4658 N$34659 N$34660 N$18116 N$18118 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4659 N$34661 N$34662 N$18120 N$18122 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4660 N$34663 N$34664 N$18124 N$18126 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4661 N$34665 N$34666 N$18128 N$18130 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4662 N$34667 N$34668 N$18132 N$18134 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4663 N$34669 N$34670 N$18136 N$18138 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4664 N$34671 N$34672 N$18140 N$18142 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4665 N$34673 N$34674 N$18144 N$18146 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4666 N$34675 N$34676 N$18148 N$18150 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4667 N$34677 N$34678 N$18152 N$18154 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4668 N$34679 N$34680 N$18156 N$18158 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4669 N$34681 N$34682 N$18160 N$18162 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4670 N$34683 N$34684 N$18164 N$18166 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4671 N$34685 N$34686 N$18168 N$18170 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4672 N$34687 N$34688 N$18172 N$26239 BDC_switch_ideal library="Design kits/capstone" sch_x=-254 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4673 N$17921 N$17923 N$25985 N$18174 "Waveguide Crossing" sch_x=-252 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4674 N$17925 N$17927 N$18176 N$18178 "Waveguide Crossing" sch_x=-252 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4675 N$17929 N$17931 N$18180 N$18182 "Waveguide Crossing" sch_x=-252 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4676 N$17933 N$17935 N$18184 N$18186 "Waveguide Crossing" sch_x=-252 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4677 N$17937 N$17939 N$18188 N$18190 "Waveguide Crossing" sch_x=-252 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4678 N$17941 N$17943 N$18192 N$18194 "Waveguide Crossing" sch_x=-252 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4679 N$17945 N$17947 N$18196 N$18198 "Waveguide Crossing" sch_x=-252 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4680 N$17949 N$17951 N$18200 N$18202 "Waveguide Crossing" sch_x=-252 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4681 N$17953 N$17955 N$18204 N$18206 "Waveguide Crossing" sch_x=-252 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4682 N$17957 N$17959 N$18208 N$18210 "Waveguide Crossing" sch_x=-252 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4683 N$17961 N$17963 N$18212 N$18214 "Waveguide Crossing" sch_x=-252 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4684 N$17965 N$17967 N$18216 N$18218 "Waveguide Crossing" sch_x=-252 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4685 N$17969 N$17971 N$18220 N$18222 "Waveguide Crossing" sch_x=-252 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4686 N$17973 N$17975 N$18224 N$18226 "Waveguide Crossing" sch_x=-252 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4687 N$17977 N$17979 N$18228 N$18230 "Waveguide Crossing" sch_x=-252 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4688 N$17981 N$17983 N$18232 N$18234 "Waveguide Crossing" sch_x=-252 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4689 N$17985 N$17987 N$18236 N$18238 "Waveguide Crossing" sch_x=-252 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4690 N$17989 N$17991 N$18240 N$18242 "Waveguide Crossing" sch_x=-252 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4691 N$17993 N$17995 N$18244 N$18246 "Waveguide Crossing" sch_x=-252 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4692 N$17997 N$17999 N$18248 N$18250 "Waveguide Crossing" sch_x=-252 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4693 N$18001 N$18003 N$18252 N$18254 "Waveguide Crossing" sch_x=-252 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4694 N$18005 N$18007 N$18256 N$18258 "Waveguide Crossing" sch_x=-252 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4695 N$18009 N$18011 N$18260 N$18262 "Waveguide Crossing" sch_x=-252 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4696 N$18013 N$18015 N$18264 N$18266 "Waveguide Crossing" sch_x=-252 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4697 N$18017 N$18019 N$18268 N$18270 "Waveguide Crossing" sch_x=-252 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4698 N$18021 N$18023 N$18272 N$18274 "Waveguide Crossing" sch_x=-252 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4699 N$18025 N$18027 N$18276 N$18278 "Waveguide Crossing" sch_x=-252 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4700 N$18029 N$18031 N$18280 N$18282 "Waveguide Crossing" sch_x=-252 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4701 N$18033 N$18035 N$18284 N$18286 "Waveguide Crossing" sch_x=-252 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4702 N$18037 N$18039 N$18288 N$18290 "Waveguide Crossing" sch_x=-252 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4703 N$18041 N$18043 N$18292 N$18294 "Waveguide Crossing" sch_x=-252 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4704 N$18045 N$18047 N$18296 N$18298 "Waveguide Crossing" sch_x=-252 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4705 N$18049 N$18051 N$18300 N$18302 "Waveguide Crossing" sch_x=-252 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4706 N$18053 N$18055 N$18304 N$18306 "Waveguide Crossing" sch_x=-252 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4707 N$18057 N$18059 N$18308 N$18310 "Waveguide Crossing" sch_x=-252 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4708 N$18061 N$18063 N$18312 N$18314 "Waveguide Crossing" sch_x=-252 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4709 N$18065 N$18067 N$18316 N$18318 "Waveguide Crossing" sch_x=-252 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4710 N$18069 N$18071 N$18320 N$18322 "Waveguide Crossing" sch_x=-252 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4711 N$18073 N$18075 N$18324 N$18326 "Waveguide Crossing" sch_x=-252 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4712 N$18077 N$18079 N$18328 N$18330 "Waveguide Crossing" sch_x=-252 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4713 N$18081 N$18083 N$18332 N$18334 "Waveguide Crossing" sch_x=-252 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4714 N$18085 N$18087 N$18336 N$18338 "Waveguide Crossing" sch_x=-252 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4715 N$18089 N$18091 N$18340 N$18342 "Waveguide Crossing" sch_x=-252 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4716 N$18093 N$18095 N$18344 N$18346 "Waveguide Crossing" sch_x=-252 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4717 N$18097 N$18099 N$18348 N$18350 "Waveguide Crossing" sch_x=-252 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4718 N$18101 N$18103 N$18352 N$18354 "Waveguide Crossing" sch_x=-252 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4719 N$18105 N$18107 N$18356 N$18358 "Waveguide Crossing" sch_x=-252 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4720 N$18109 N$18111 N$18360 N$18362 "Waveguide Crossing" sch_x=-252 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4721 N$18113 N$18115 N$18364 N$18366 "Waveguide Crossing" sch_x=-252 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4722 N$18117 N$18119 N$18368 N$18370 "Waveguide Crossing" sch_x=-252 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4723 N$18121 N$18123 N$18372 N$18374 "Waveguide Crossing" sch_x=-252 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4724 N$18125 N$18127 N$18376 N$18378 "Waveguide Crossing" sch_x=-252 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4725 N$18129 N$18131 N$18380 N$18382 "Waveguide Crossing" sch_x=-252 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4726 N$18133 N$18135 N$18384 N$18386 "Waveguide Crossing" sch_x=-252 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4727 N$18137 N$18139 N$18388 N$18390 "Waveguide Crossing" sch_x=-252 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4728 N$18141 N$18143 N$18392 N$18394 "Waveguide Crossing" sch_x=-252 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4729 N$18145 N$18147 N$18396 N$18398 "Waveguide Crossing" sch_x=-252 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4730 N$18149 N$18151 N$18400 N$18402 "Waveguide Crossing" sch_x=-252 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4731 N$18153 N$18155 N$18404 N$18406 "Waveguide Crossing" sch_x=-252 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4732 N$18157 N$18159 N$18408 N$18410 "Waveguide Crossing" sch_x=-252 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4733 N$18161 N$18163 N$18412 N$18414 "Waveguide Crossing" sch_x=-252 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4734 N$18165 N$18167 N$18416 N$18418 "Waveguide Crossing" sch_x=-252 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4735 N$18169 N$18171 N$18420 N$26235 "Waveguide Crossing" sch_x=-252 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4736 N$18173 N$18175 N$25987 N$18422 "Waveguide Crossing" sch_x=-250 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4737 N$18177 N$18179 N$18424 N$18426 "Waveguide Crossing" sch_x=-250 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4738 N$18181 N$18183 N$18428 N$18430 "Waveguide Crossing" sch_x=-250 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4739 N$18185 N$18187 N$18432 N$18434 "Waveguide Crossing" sch_x=-250 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4740 N$18189 N$18191 N$18436 N$18438 "Waveguide Crossing" sch_x=-250 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4741 N$18193 N$18195 N$18440 N$18442 "Waveguide Crossing" sch_x=-250 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4742 N$18197 N$18199 N$18444 N$18446 "Waveguide Crossing" sch_x=-250 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4743 N$18201 N$18203 N$18448 N$18450 "Waveguide Crossing" sch_x=-250 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4744 N$18205 N$18207 N$18452 N$18454 "Waveguide Crossing" sch_x=-250 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4745 N$18209 N$18211 N$18456 N$18458 "Waveguide Crossing" sch_x=-250 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4746 N$18213 N$18215 N$18460 N$18462 "Waveguide Crossing" sch_x=-250 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4747 N$18217 N$18219 N$18464 N$18466 "Waveguide Crossing" sch_x=-250 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4748 N$18221 N$18223 N$18468 N$18470 "Waveguide Crossing" sch_x=-250 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4749 N$18225 N$18227 N$18472 N$18474 "Waveguide Crossing" sch_x=-250 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4750 N$18229 N$18231 N$18476 N$18478 "Waveguide Crossing" sch_x=-250 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4751 N$18233 N$18235 N$18480 N$18482 "Waveguide Crossing" sch_x=-250 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4752 N$18237 N$18239 N$18484 N$18486 "Waveguide Crossing" sch_x=-250 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4753 N$18241 N$18243 N$18488 N$18490 "Waveguide Crossing" sch_x=-250 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4754 N$18245 N$18247 N$18492 N$18494 "Waveguide Crossing" sch_x=-250 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4755 N$18249 N$18251 N$18496 N$18498 "Waveguide Crossing" sch_x=-250 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4756 N$18253 N$18255 N$18500 N$18502 "Waveguide Crossing" sch_x=-250 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4757 N$18257 N$18259 N$18504 N$18506 "Waveguide Crossing" sch_x=-250 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4758 N$18261 N$18263 N$18508 N$18510 "Waveguide Crossing" sch_x=-250 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4759 N$18265 N$18267 N$18512 N$18514 "Waveguide Crossing" sch_x=-250 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4760 N$18269 N$18271 N$18516 N$18518 "Waveguide Crossing" sch_x=-250 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4761 N$18273 N$18275 N$18520 N$18522 "Waveguide Crossing" sch_x=-250 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4762 N$18277 N$18279 N$18524 N$18526 "Waveguide Crossing" sch_x=-250 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4763 N$18281 N$18283 N$18528 N$18530 "Waveguide Crossing" sch_x=-250 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4764 N$18285 N$18287 N$18532 N$18534 "Waveguide Crossing" sch_x=-250 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4765 N$18289 N$18291 N$18536 N$18538 "Waveguide Crossing" sch_x=-250 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4766 N$18293 N$18295 N$18540 N$18542 "Waveguide Crossing" sch_x=-250 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4767 N$18297 N$18299 N$18544 N$18546 "Waveguide Crossing" sch_x=-250 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4768 N$18301 N$18303 N$18548 N$18550 "Waveguide Crossing" sch_x=-250 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4769 N$18305 N$18307 N$18552 N$18554 "Waveguide Crossing" sch_x=-250 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4770 N$18309 N$18311 N$18556 N$18558 "Waveguide Crossing" sch_x=-250 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4771 N$18313 N$18315 N$18560 N$18562 "Waveguide Crossing" sch_x=-250 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4772 N$18317 N$18319 N$18564 N$18566 "Waveguide Crossing" sch_x=-250 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4773 N$18321 N$18323 N$18568 N$18570 "Waveguide Crossing" sch_x=-250 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4774 N$18325 N$18327 N$18572 N$18574 "Waveguide Crossing" sch_x=-250 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4775 N$18329 N$18331 N$18576 N$18578 "Waveguide Crossing" sch_x=-250 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4776 N$18333 N$18335 N$18580 N$18582 "Waveguide Crossing" sch_x=-250 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4777 N$18337 N$18339 N$18584 N$18586 "Waveguide Crossing" sch_x=-250 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4778 N$18341 N$18343 N$18588 N$18590 "Waveguide Crossing" sch_x=-250 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4779 N$18345 N$18347 N$18592 N$18594 "Waveguide Crossing" sch_x=-250 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4780 N$18349 N$18351 N$18596 N$18598 "Waveguide Crossing" sch_x=-250 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4781 N$18353 N$18355 N$18600 N$18602 "Waveguide Crossing" sch_x=-250 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4782 N$18357 N$18359 N$18604 N$18606 "Waveguide Crossing" sch_x=-250 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4783 N$18361 N$18363 N$18608 N$18610 "Waveguide Crossing" sch_x=-250 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4784 N$18365 N$18367 N$18612 N$18614 "Waveguide Crossing" sch_x=-250 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4785 N$18369 N$18371 N$18616 N$18618 "Waveguide Crossing" sch_x=-250 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4786 N$18373 N$18375 N$18620 N$18622 "Waveguide Crossing" sch_x=-250 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4787 N$18377 N$18379 N$18624 N$18626 "Waveguide Crossing" sch_x=-250 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4788 N$18381 N$18383 N$18628 N$18630 "Waveguide Crossing" sch_x=-250 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4789 N$18385 N$18387 N$18632 N$18634 "Waveguide Crossing" sch_x=-250 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4790 N$18389 N$18391 N$18636 N$18638 "Waveguide Crossing" sch_x=-250 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4791 N$18393 N$18395 N$18640 N$18642 "Waveguide Crossing" sch_x=-250 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4792 N$18397 N$18399 N$18644 N$18646 "Waveguide Crossing" sch_x=-250 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4793 N$18401 N$18403 N$18648 N$18650 "Waveguide Crossing" sch_x=-250 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4794 N$18405 N$18407 N$18652 N$18654 "Waveguide Crossing" sch_x=-250 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4795 N$18409 N$18411 N$18656 N$18658 "Waveguide Crossing" sch_x=-250 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4796 N$18413 N$18415 N$18660 N$18662 "Waveguide Crossing" sch_x=-250 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4797 N$18417 N$18419 N$18664 N$26233 "Waveguide Crossing" sch_x=-250 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4798 N$18421 N$18423 N$25989 N$18666 "Waveguide Crossing" sch_x=-248 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4799 N$18425 N$18427 N$18668 N$18670 "Waveguide Crossing" sch_x=-248 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4800 N$18429 N$18431 N$18672 N$18674 "Waveguide Crossing" sch_x=-248 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4801 N$18433 N$18435 N$18676 N$18678 "Waveguide Crossing" sch_x=-248 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4802 N$18437 N$18439 N$18680 N$18682 "Waveguide Crossing" sch_x=-248 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4803 N$18441 N$18443 N$18684 N$18686 "Waveguide Crossing" sch_x=-248 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4804 N$18445 N$18447 N$18688 N$18690 "Waveguide Crossing" sch_x=-248 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4805 N$18449 N$18451 N$18692 N$18694 "Waveguide Crossing" sch_x=-248 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4806 N$18453 N$18455 N$18696 N$18698 "Waveguide Crossing" sch_x=-248 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4807 N$18457 N$18459 N$18700 N$18702 "Waveguide Crossing" sch_x=-248 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4808 N$18461 N$18463 N$18704 N$18706 "Waveguide Crossing" sch_x=-248 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4809 N$18465 N$18467 N$18708 N$18710 "Waveguide Crossing" sch_x=-248 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4810 N$18469 N$18471 N$18712 N$18714 "Waveguide Crossing" sch_x=-248 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4811 N$18473 N$18475 N$18716 N$18718 "Waveguide Crossing" sch_x=-248 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4812 N$18477 N$18479 N$18720 N$18722 "Waveguide Crossing" sch_x=-248 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4813 N$18481 N$18483 N$18724 N$18726 "Waveguide Crossing" sch_x=-248 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4814 N$18485 N$18487 N$18728 N$18730 "Waveguide Crossing" sch_x=-248 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4815 N$18489 N$18491 N$18732 N$18734 "Waveguide Crossing" sch_x=-248 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4816 N$18493 N$18495 N$18736 N$18738 "Waveguide Crossing" sch_x=-248 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4817 N$18497 N$18499 N$18740 N$18742 "Waveguide Crossing" sch_x=-248 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4818 N$18501 N$18503 N$18744 N$18746 "Waveguide Crossing" sch_x=-248 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4819 N$18505 N$18507 N$18748 N$18750 "Waveguide Crossing" sch_x=-248 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4820 N$18509 N$18511 N$18752 N$18754 "Waveguide Crossing" sch_x=-248 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4821 N$18513 N$18515 N$18756 N$18758 "Waveguide Crossing" sch_x=-248 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4822 N$18517 N$18519 N$18760 N$18762 "Waveguide Crossing" sch_x=-248 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4823 N$18521 N$18523 N$18764 N$18766 "Waveguide Crossing" sch_x=-248 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4824 N$18525 N$18527 N$18768 N$18770 "Waveguide Crossing" sch_x=-248 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4825 N$18529 N$18531 N$18772 N$18774 "Waveguide Crossing" sch_x=-248 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4826 N$18533 N$18535 N$18776 N$18778 "Waveguide Crossing" sch_x=-248 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4827 N$18537 N$18539 N$18780 N$18782 "Waveguide Crossing" sch_x=-248 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4828 N$18541 N$18543 N$18784 N$18786 "Waveguide Crossing" sch_x=-248 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4829 N$18545 N$18547 N$18788 N$18790 "Waveguide Crossing" sch_x=-248 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4830 N$18549 N$18551 N$18792 N$18794 "Waveguide Crossing" sch_x=-248 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4831 N$18553 N$18555 N$18796 N$18798 "Waveguide Crossing" sch_x=-248 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4832 N$18557 N$18559 N$18800 N$18802 "Waveguide Crossing" sch_x=-248 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4833 N$18561 N$18563 N$18804 N$18806 "Waveguide Crossing" sch_x=-248 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4834 N$18565 N$18567 N$18808 N$18810 "Waveguide Crossing" sch_x=-248 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4835 N$18569 N$18571 N$18812 N$18814 "Waveguide Crossing" sch_x=-248 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4836 N$18573 N$18575 N$18816 N$18818 "Waveguide Crossing" sch_x=-248 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4837 N$18577 N$18579 N$18820 N$18822 "Waveguide Crossing" sch_x=-248 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4838 N$18581 N$18583 N$18824 N$18826 "Waveguide Crossing" sch_x=-248 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4839 N$18585 N$18587 N$18828 N$18830 "Waveguide Crossing" sch_x=-248 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4840 N$18589 N$18591 N$18832 N$18834 "Waveguide Crossing" sch_x=-248 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4841 N$18593 N$18595 N$18836 N$18838 "Waveguide Crossing" sch_x=-248 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4842 N$18597 N$18599 N$18840 N$18842 "Waveguide Crossing" sch_x=-248 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4843 N$18601 N$18603 N$18844 N$18846 "Waveguide Crossing" sch_x=-248 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4844 N$18605 N$18607 N$18848 N$18850 "Waveguide Crossing" sch_x=-248 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4845 N$18609 N$18611 N$18852 N$18854 "Waveguide Crossing" sch_x=-248 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4846 N$18613 N$18615 N$18856 N$18858 "Waveguide Crossing" sch_x=-248 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4847 N$18617 N$18619 N$18860 N$18862 "Waveguide Crossing" sch_x=-248 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4848 N$18621 N$18623 N$18864 N$18866 "Waveguide Crossing" sch_x=-248 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4849 N$18625 N$18627 N$18868 N$18870 "Waveguide Crossing" sch_x=-248 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4850 N$18629 N$18631 N$18872 N$18874 "Waveguide Crossing" sch_x=-248 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4851 N$18633 N$18635 N$18876 N$18878 "Waveguide Crossing" sch_x=-248 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4852 N$18637 N$18639 N$18880 N$18882 "Waveguide Crossing" sch_x=-248 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4853 N$18641 N$18643 N$18884 N$18886 "Waveguide Crossing" sch_x=-248 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4854 N$18645 N$18647 N$18888 N$18890 "Waveguide Crossing" sch_x=-248 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4855 N$18649 N$18651 N$18892 N$18894 "Waveguide Crossing" sch_x=-248 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4856 N$18653 N$18655 N$18896 N$18898 "Waveguide Crossing" sch_x=-248 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4857 N$18657 N$18659 N$18900 N$18902 "Waveguide Crossing" sch_x=-248 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4858 N$18661 N$18663 N$18904 N$26231 "Waveguide Crossing" sch_x=-248 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4859 N$18665 N$18667 N$25991 N$18906 "Waveguide Crossing" sch_x=-246 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4860 N$18669 N$18671 N$18908 N$18910 "Waveguide Crossing" sch_x=-246 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4861 N$18673 N$18675 N$18912 N$18914 "Waveguide Crossing" sch_x=-246 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4862 N$18677 N$18679 N$18916 N$18918 "Waveguide Crossing" sch_x=-246 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4863 N$18681 N$18683 N$18920 N$18922 "Waveguide Crossing" sch_x=-246 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4864 N$18685 N$18687 N$18924 N$18926 "Waveguide Crossing" sch_x=-246 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4865 N$18689 N$18691 N$18928 N$18930 "Waveguide Crossing" sch_x=-246 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4866 N$18693 N$18695 N$18932 N$18934 "Waveguide Crossing" sch_x=-246 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4867 N$18697 N$18699 N$18936 N$18938 "Waveguide Crossing" sch_x=-246 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4868 N$18701 N$18703 N$18940 N$18942 "Waveguide Crossing" sch_x=-246 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4869 N$18705 N$18707 N$18944 N$18946 "Waveguide Crossing" sch_x=-246 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4870 N$18709 N$18711 N$18948 N$18950 "Waveguide Crossing" sch_x=-246 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4871 N$18713 N$18715 N$18952 N$18954 "Waveguide Crossing" sch_x=-246 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4872 N$18717 N$18719 N$18956 N$18958 "Waveguide Crossing" sch_x=-246 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4873 N$18721 N$18723 N$18960 N$18962 "Waveguide Crossing" sch_x=-246 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4874 N$18725 N$18727 N$18964 N$18966 "Waveguide Crossing" sch_x=-246 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4875 N$18729 N$18731 N$18968 N$18970 "Waveguide Crossing" sch_x=-246 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4876 N$18733 N$18735 N$18972 N$18974 "Waveguide Crossing" sch_x=-246 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4877 N$18737 N$18739 N$18976 N$18978 "Waveguide Crossing" sch_x=-246 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4878 N$18741 N$18743 N$18980 N$18982 "Waveguide Crossing" sch_x=-246 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4879 N$18745 N$18747 N$18984 N$18986 "Waveguide Crossing" sch_x=-246 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4880 N$18749 N$18751 N$18988 N$18990 "Waveguide Crossing" sch_x=-246 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4881 N$18753 N$18755 N$18992 N$18994 "Waveguide Crossing" sch_x=-246 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4882 N$18757 N$18759 N$18996 N$18998 "Waveguide Crossing" sch_x=-246 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4883 N$18761 N$18763 N$19000 N$19002 "Waveguide Crossing" sch_x=-246 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4884 N$18765 N$18767 N$19004 N$19006 "Waveguide Crossing" sch_x=-246 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4885 N$18769 N$18771 N$19008 N$19010 "Waveguide Crossing" sch_x=-246 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4886 N$18773 N$18775 N$19012 N$19014 "Waveguide Crossing" sch_x=-246 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4887 N$18777 N$18779 N$19016 N$19018 "Waveguide Crossing" sch_x=-246 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4888 N$18781 N$18783 N$19020 N$19022 "Waveguide Crossing" sch_x=-246 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4889 N$18785 N$18787 N$19024 N$19026 "Waveguide Crossing" sch_x=-246 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4890 N$18789 N$18791 N$19028 N$19030 "Waveguide Crossing" sch_x=-246 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4891 N$18793 N$18795 N$19032 N$19034 "Waveguide Crossing" sch_x=-246 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4892 N$18797 N$18799 N$19036 N$19038 "Waveguide Crossing" sch_x=-246 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4893 N$18801 N$18803 N$19040 N$19042 "Waveguide Crossing" sch_x=-246 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4894 N$18805 N$18807 N$19044 N$19046 "Waveguide Crossing" sch_x=-246 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4895 N$18809 N$18811 N$19048 N$19050 "Waveguide Crossing" sch_x=-246 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4896 N$18813 N$18815 N$19052 N$19054 "Waveguide Crossing" sch_x=-246 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4897 N$18817 N$18819 N$19056 N$19058 "Waveguide Crossing" sch_x=-246 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4898 N$18821 N$18823 N$19060 N$19062 "Waveguide Crossing" sch_x=-246 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4899 N$18825 N$18827 N$19064 N$19066 "Waveguide Crossing" sch_x=-246 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4900 N$18829 N$18831 N$19068 N$19070 "Waveguide Crossing" sch_x=-246 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4901 N$18833 N$18835 N$19072 N$19074 "Waveguide Crossing" sch_x=-246 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4902 N$18837 N$18839 N$19076 N$19078 "Waveguide Crossing" sch_x=-246 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4903 N$18841 N$18843 N$19080 N$19082 "Waveguide Crossing" sch_x=-246 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4904 N$18845 N$18847 N$19084 N$19086 "Waveguide Crossing" sch_x=-246 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4905 N$18849 N$18851 N$19088 N$19090 "Waveguide Crossing" sch_x=-246 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4906 N$18853 N$18855 N$19092 N$19094 "Waveguide Crossing" sch_x=-246 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4907 N$18857 N$18859 N$19096 N$19098 "Waveguide Crossing" sch_x=-246 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4908 N$18861 N$18863 N$19100 N$19102 "Waveguide Crossing" sch_x=-246 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4909 N$18865 N$18867 N$19104 N$19106 "Waveguide Crossing" sch_x=-246 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4910 N$18869 N$18871 N$19108 N$19110 "Waveguide Crossing" sch_x=-246 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4911 N$18873 N$18875 N$19112 N$19114 "Waveguide Crossing" sch_x=-246 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4912 N$18877 N$18879 N$19116 N$19118 "Waveguide Crossing" sch_x=-246 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4913 N$18881 N$18883 N$19120 N$19122 "Waveguide Crossing" sch_x=-246 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4914 N$18885 N$18887 N$19124 N$19126 "Waveguide Crossing" sch_x=-246 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4915 N$18889 N$18891 N$19128 N$19130 "Waveguide Crossing" sch_x=-246 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4916 N$18893 N$18895 N$19132 N$19134 "Waveguide Crossing" sch_x=-246 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4917 N$18897 N$18899 N$19136 N$19138 "Waveguide Crossing" sch_x=-246 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4918 N$18901 N$18903 N$19140 N$26229 "Waveguide Crossing" sch_x=-246 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4919 N$18905 N$18907 N$25993 N$19142 "Waveguide Crossing" sch_x=-244 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4920 N$18909 N$18911 N$19144 N$19146 "Waveguide Crossing" sch_x=-244 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4921 N$18913 N$18915 N$19148 N$19150 "Waveguide Crossing" sch_x=-244 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4922 N$18917 N$18919 N$19152 N$19154 "Waveguide Crossing" sch_x=-244 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4923 N$18921 N$18923 N$19156 N$19158 "Waveguide Crossing" sch_x=-244 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4924 N$18925 N$18927 N$19160 N$19162 "Waveguide Crossing" sch_x=-244 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4925 N$18929 N$18931 N$19164 N$19166 "Waveguide Crossing" sch_x=-244 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4926 N$18933 N$18935 N$19168 N$19170 "Waveguide Crossing" sch_x=-244 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4927 N$18937 N$18939 N$19172 N$19174 "Waveguide Crossing" sch_x=-244 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4928 N$18941 N$18943 N$19176 N$19178 "Waveguide Crossing" sch_x=-244 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4929 N$18945 N$18947 N$19180 N$19182 "Waveguide Crossing" sch_x=-244 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4930 N$18949 N$18951 N$19184 N$19186 "Waveguide Crossing" sch_x=-244 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4931 N$18953 N$18955 N$19188 N$19190 "Waveguide Crossing" sch_x=-244 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4932 N$18957 N$18959 N$19192 N$19194 "Waveguide Crossing" sch_x=-244 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4933 N$18961 N$18963 N$19196 N$19198 "Waveguide Crossing" sch_x=-244 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4934 N$18965 N$18967 N$19200 N$19202 "Waveguide Crossing" sch_x=-244 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4935 N$18969 N$18971 N$19204 N$19206 "Waveguide Crossing" sch_x=-244 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4936 N$18973 N$18975 N$19208 N$19210 "Waveguide Crossing" sch_x=-244 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4937 N$18977 N$18979 N$19212 N$19214 "Waveguide Crossing" sch_x=-244 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4938 N$18981 N$18983 N$19216 N$19218 "Waveguide Crossing" sch_x=-244 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4939 N$18985 N$18987 N$19220 N$19222 "Waveguide Crossing" sch_x=-244 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4940 N$18989 N$18991 N$19224 N$19226 "Waveguide Crossing" sch_x=-244 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4941 N$18993 N$18995 N$19228 N$19230 "Waveguide Crossing" sch_x=-244 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4942 N$18997 N$18999 N$19232 N$19234 "Waveguide Crossing" sch_x=-244 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4943 N$19001 N$19003 N$19236 N$19238 "Waveguide Crossing" sch_x=-244 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4944 N$19005 N$19007 N$19240 N$19242 "Waveguide Crossing" sch_x=-244 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4945 N$19009 N$19011 N$19244 N$19246 "Waveguide Crossing" sch_x=-244 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4946 N$19013 N$19015 N$19248 N$19250 "Waveguide Crossing" sch_x=-244 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4947 N$19017 N$19019 N$19252 N$19254 "Waveguide Crossing" sch_x=-244 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4948 N$19021 N$19023 N$19256 N$19258 "Waveguide Crossing" sch_x=-244 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4949 N$19025 N$19027 N$19260 N$19262 "Waveguide Crossing" sch_x=-244 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4950 N$19029 N$19031 N$19264 N$19266 "Waveguide Crossing" sch_x=-244 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4951 N$19033 N$19035 N$19268 N$19270 "Waveguide Crossing" sch_x=-244 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4952 N$19037 N$19039 N$19272 N$19274 "Waveguide Crossing" sch_x=-244 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4953 N$19041 N$19043 N$19276 N$19278 "Waveguide Crossing" sch_x=-244 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4954 N$19045 N$19047 N$19280 N$19282 "Waveguide Crossing" sch_x=-244 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4955 N$19049 N$19051 N$19284 N$19286 "Waveguide Crossing" sch_x=-244 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4956 N$19053 N$19055 N$19288 N$19290 "Waveguide Crossing" sch_x=-244 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4957 N$19057 N$19059 N$19292 N$19294 "Waveguide Crossing" sch_x=-244 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4958 N$19061 N$19063 N$19296 N$19298 "Waveguide Crossing" sch_x=-244 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4959 N$19065 N$19067 N$19300 N$19302 "Waveguide Crossing" sch_x=-244 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4960 N$19069 N$19071 N$19304 N$19306 "Waveguide Crossing" sch_x=-244 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4961 N$19073 N$19075 N$19308 N$19310 "Waveguide Crossing" sch_x=-244 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4962 N$19077 N$19079 N$19312 N$19314 "Waveguide Crossing" sch_x=-244 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4963 N$19081 N$19083 N$19316 N$19318 "Waveguide Crossing" sch_x=-244 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4964 N$19085 N$19087 N$19320 N$19322 "Waveguide Crossing" sch_x=-244 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4965 N$19089 N$19091 N$19324 N$19326 "Waveguide Crossing" sch_x=-244 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4966 N$19093 N$19095 N$19328 N$19330 "Waveguide Crossing" sch_x=-244 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4967 N$19097 N$19099 N$19332 N$19334 "Waveguide Crossing" sch_x=-244 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4968 N$19101 N$19103 N$19336 N$19338 "Waveguide Crossing" sch_x=-244 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4969 N$19105 N$19107 N$19340 N$19342 "Waveguide Crossing" sch_x=-244 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4970 N$19109 N$19111 N$19344 N$19346 "Waveguide Crossing" sch_x=-244 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4971 N$19113 N$19115 N$19348 N$19350 "Waveguide Crossing" sch_x=-244 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4972 N$19117 N$19119 N$19352 N$19354 "Waveguide Crossing" sch_x=-244 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4973 N$19121 N$19123 N$19356 N$19358 "Waveguide Crossing" sch_x=-244 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4974 N$19125 N$19127 N$19360 N$19362 "Waveguide Crossing" sch_x=-244 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4975 N$19129 N$19131 N$19364 N$19366 "Waveguide Crossing" sch_x=-244 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4976 N$19133 N$19135 N$19368 N$19370 "Waveguide Crossing" sch_x=-244 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4977 N$19137 N$19139 N$19372 N$26227 "Waveguide Crossing" sch_x=-244 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4978 N$19141 N$19143 N$25995 N$19374 "Waveguide Crossing" sch_x=-242 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4979 N$19145 N$19147 N$19376 N$19378 "Waveguide Crossing" sch_x=-242 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4980 N$19149 N$19151 N$19380 N$19382 "Waveguide Crossing" sch_x=-242 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4981 N$19153 N$19155 N$19384 N$19386 "Waveguide Crossing" sch_x=-242 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4982 N$19157 N$19159 N$19388 N$19390 "Waveguide Crossing" sch_x=-242 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4983 N$19161 N$19163 N$19392 N$19394 "Waveguide Crossing" sch_x=-242 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4984 N$19165 N$19167 N$19396 N$19398 "Waveguide Crossing" sch_x=-242 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4985 N$19169 N$19171 N$19400 N$19402 "Waveguide Crossing" sch_x=-242 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4986 N$19173 N$19175 N$19404 N$19406 "Waveguide Crossing" sch_x=-242 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4987 N$19177 N$19179 N$19408 N$19410 "Waveguide Crossing" sch_x=-242 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4988 N$19181 N$19183 N$19412 N$19414 "Waveguide Crossing" sch_x=-242 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4989 N$19185 N$19187 N$19416 N$19418 "Waveguide Crossing" sch_x=-242 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4990 N$19189 N$19191 N$19420 N$19422 "Waveguide Crossing" sch_x=-242 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4991 N$19193 N$19195 N$19424 N$19426 "Waveguide Crossing" sch_x=-242 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4992 N$19197 N$19199 N$19428 N$19430 "Waveguide Crossing" sch_x=-242 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4993 N$19201 N$19203 N$19432 N$19434 "Waveguide Crossing" sch_x=-242 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4994 N$19205 N$19207 N$19436 N$19438 "Waveguide Crossing" sch_x=-242 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4995 N$19209 N$19211 N$19440 N$19442 "Waveguide Crossing" sch_x=-242 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4996 N$19213 N$19215 N$19444 N$19446 "Waveguide Crossing" sch_x=-242 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4997 N$19217 N$19219 N$19448 N$19450 "Waveguide Crossing" sch_x=-242 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4998 N$19221 N$19223 N$19452 N$19454 "Waveguide Crossing" sch_x=-242 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4999 N$19225 N$19227 N$19456 N$19458 "Waveguide Crossing" sch_x=-242 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5000 N$19229 N$19231 N$19460 N$19462 "Waveguide Crossing" sch_x=-242 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5001 N$19233 N$19235 N$19464 N$19466 "Waveguide Crossing" sch_x=-242 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5002 N$19237 N$19239 N$19468 N$19470 "Waveguide Crossing" sch_x=-242 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5003 N$19241 N$19243 N$19472 N$19474 "Waveguide Crossing" sch_x=-242 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5004 N$19245 N$19247 N$19476 N$19478 "Waveguide Crossing" sch_x=-242 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5005 N$19249 N$19251 N$19480 N$19482 "Waveguide Crossing" sch_x=-242 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5006 N$19253 N$19255 N$19484 N$19486 "Waveguide Crossing" sch_x=-242 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5007 N$19257 N$19259 N$19488 N$19490 "Waveguide Crossing" sch_x=-242 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5008 N$19261 N$19263 N$19492 N$19494 "Waveguide Crossing" sch_x=-242 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5009 N$19265 N$19267 N$19496 N$19498 "Waveguide Crossing" sch_x=-242 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5010 N$19269 N$19271 N$19500 N$19502 "Waveguide Crossing" sch_x=-242 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5011 N$19273 N$19275 N$19504 N$19506 "Waveguide Crossing" sch_x=-242 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5012 N$19277 N$19279 N$19508 N$19510 "Waveguide Crossing" sch_x=-242 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5013 N$19281 N$19283 N$19512 N$19514 "Waveguide Crossing" sch_x=-242 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5014 N$19285 N$19287 N$19516 N$19518 "Waveguide Crossing" sch_x=-242 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5015 N$19289 N$19291 N$19520 N$19522 "Waveguide Crossing" sch_x=-242 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5016 N$19293 N$19295 N$19524 N$19526 "Waveguide Crossing" sch_x=-242 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5017 N$19297 N$19299 N$19528 N$19530 "Waveguide Crossing" sch_x=-242 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5018 N$19301 N$19303 N$19532 N$19534 "Waveguide Crossing" sch_x=-242 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5019 N$19305 N$19307 N$19536 N$19538 "Waveguide Crossing" sch_x=-242 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5020 N$19309 N$19311 N$19540 N$19542 "Waveguide Crossing" sch_x=-242 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5021 N$19313 N$19315 N$19544 N$19546 "Waveguide Crossing" sch_x=-242 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5022 N$19317 N$19319 N$19548 N$19550 "Waveguide Crossing" sch_x=-242 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5023 N$19321 N$19323 N$19552 N$19554 "Waveguide Crossing" sch_x=-242 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5024 N$19325 N$19327 N$19556 N$19558 "Waveguide Crossing" sch_x=-242 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5025 N$19329 N$19331 N$19560 N$19562 "Waveguide Crossing" sch_x=-242 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5026 N$19333 N$19335 N$19564 N$19566 "Waveguide Crossing" sch_x=-242 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5027 N$19337 N$19339 N$19568 N$19570 "Waveguide Crossing" sch_x=-242 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5028 N$19341 N$19343 N$19572 N$19574 "Waveguide Crossing" sch_x=-242 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5029 N$19345 N$19347 N$19576 N$19578 "Waveguide Crossing" sch_x=-242 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5030 N$19349 N$19351 N$19580 N$19582 "Waveguide Crossing" sch_x=-242 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5031 N$19353 N$19355 N$19584 N$19586 "Waveguide Crossing" sch_x=-242 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5032 N$19357 N$19359 N$19588 N$19590 "Waveguide Crossing" sch_x=-242 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5033 N$19361 N$19363 N$19592 N$19594 "Waveguide Crossing" sch_x=-242 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5034 N$19365 N$19367 N$19596 N$19598 "Waveguide Crossing" sch_x=-242 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5035 N$19369 N$19371 N$19600 N$26225 "Waveguide Crossing" sch_x=-242 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5036 N$19373 N$19375 N$25997 N$19602 "Waveguide Crossing" sch_x=-240 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5037 N$19377 N$19379 N$19604 N$19606 "Waveguide Crossing" sch_x=-240 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5038 N$19381 N$19383 N$19608 N$19610 "Waveguide Crossing" sch_x=-240 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5039 N$19385 N$19387 N$19612 N$19614 "Waveguide Crossing" sch_x=-240 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5040 N$19389 N$19391 N$19616 N$19618 "Waveguide Crossing" sch_x=-240 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5041 N$19393 N$19395 N$19620 N$19622 "Waveguide Crossing" sch_x=-240 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5042 N$19397 N$19399 N$19624 N$19626 "Waveguide Crossing" sch_x=-240 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5043 N$19401 N$19403 N$19628 N$19630 "Waveguide Crossing" sch_x=-240 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5044 N$19405 N$19407 N$19632 N$19634 "Waveguide Crossing" sch_x=-240 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5045 N$19409 N$19411 N$19636 N$19638 "Waveguide Crossing" sch_x=-240 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5046 N$19413 N$19415 N$19640 N$19642 "Waveguide Crossing" sch_x=-240 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5047 N$19417 N$19419 N$19644 N$19646 "Waveguide Crossing" sch_x=-240 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5048 N$19421 N$19423 N$19648 N$19650 "Waveguide Crossing" sch_x=-240 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5049 N$19425 N$19427 N$19652 N$19654 "Waveguide Crossing" sch_x=-240 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5050 N$19429 N$19431 N$19656 N$19658 "Waveguide Crossing" sch_x=-240 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5051 N$19433 N$19435 N$19660 N$19662 "Waveguide Crossing" sch_x=-240 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5052 N$19437 N$19439 N$19664 N$19666 "Waveguide Crossing" sch_x=-240 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5053 N$19441 N$19443 N$19668 N$19670 "Waveguide Crossing" sch_x=-240 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5054 N$19445 N$19447 N$19672 N$19674 "Waveguide Crossing" sch_x=-240 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5055 N$19449 N$19451 N$19676 N$19678 "Waveguide Crossing" sch_x=-240 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5056 N$19453 N$19455 N$19680 N$19682 "Waveguide Crossing" sch_x=-240 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5057 N$19457 N$19459 N$19684 N$19686 "Waveguide Crossing" sch_x=-240 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5058 N$19461 N$19463 N$19688 N$19690 "Waveguide Crossing" sch_x=-240 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5059 N$19465 N$19467 N$19692 N$19694 "Waveguide Crossing" sch_x=-240 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5060 N$19469 N$19471 N$19696 N$19698 "Waveguide Crossing" sch_x=-240 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5061 N$19473 N$19475 N$19700 N$19702 "Waveguide Crossing" sch_x=-240 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5062 N$19477 N$19479 N$19704 N$19706 "Waveguide Crossing" sch_x=-240 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5063 N$19481 N$19483 N$19708 N$19710 "Waveguide Crossing" sch_x=-240 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5064 N$19485 N$19487 N$19712 N$19714 "Waveguide Crossing" sch_x=-240 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5065 N$19489 N$19491 N$19716 N$19718 "Waveguide Crossing" sch_x=-240 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5066 N$19493 N$19495 N$19720 N$19722 "Waveguide Crossing" sch_x=-240 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5067 N$19497 N$19499 N$19724 N$19726 "Waveguide Crossing" sch_x=-240 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5068 N$19501 N$19503 N$19728 N$19730 "Waveguide Crossing" sch_x=-240 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5069 N$19505 N$19507 N$19732 N$19734 "Waveguide Crossing" sch_x=-240 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5070 N$19509 N$19511 N$19736 N$19738 "Waveguide Crossing" sch_x=-240 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5071 N$19513 N$19515 N$19740 N$19742 "Waveguide Crossing" sch_x=-240 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5072 N$19517 N$19519 N$19744 N$19746 "Waveguide Crossing" sch_x=-240 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5073 N$19521 N$19523 N$19748 N$19750 "Waveguide Crossing" sch_x=-240 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5074 N$19525 N$19527 N$19752 N$19754 "Waveguide Crossing" sch_x=-240 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5075 N$19529 N$19531 N$19756 N$19758 "Waveguide Crossing" sch_x=-240 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5076 N$19533 N$19535 N$19760 N$19762 "Waveguide Crossing" sch_x=-240 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5077 N$19537 N$19539 N$19764 N$19766 "Waveguide Crossing" sch_x=-240 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5078 N$19541 N$19543 N$19768 N$19770 "Waveguide Crossing" sch_x=-240 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5079 N$19545 N$19547 N$19772 N$19774 "Waveguide Crossing" sch_x=-240 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5080 N$19549 N$19551 N$19776 N$19778 "Waveguide Crossing" sch_x=-240 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5081 N$19553 N$19555 N$19780 N$19782 "Waveguide Crossing" sch_x=-240 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5082 N$19557 N$19559 N$19784 N$19786 "Waveguide Crossing" sch_x=-240 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5083 N$19561 N$19563 N$19788 N$19790 "Waveguide Crossing" sch_x=-240 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5084 N$19565 N$19567 N$19792 N$19794 "Waveguide Crossing" sch_x=-240 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5085 N$19569 N$19571 N$19796 N$19798 "Waveguide Crossing" sch_x=-240 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5086 N$19573 N$19575 N$19800 N$19802 "Waveguide Crossing" sch_x=-240 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5087 N$19577 N$19579 N$19804 N$19806 "Waveguide Crossing" sch_x=-240 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5088 N$19581 N$19583 N$19808 N$19810 "Waveguide Crossing" sch_x=-240 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5089 N$19585 N$19587 N$19812 N$19814 "Waveguide Crossing" sch_x=-240 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5090 N$19589 N$19591 N$19816 N$19818 "Waveguide Crossing" sch_x=-240 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5091 N$19593 N$19595 N$19820 N$19822 "Waveguide Crossing" sch_x=-240 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5092 N$19597 N$19599 N$19824 N$26223 "Waveguide Crossing" sch_x=-240 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5093 N$19601 N$19603 N$25999 N$19826 "Waveguide Crossing" sch_x=-238 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5094 N$19605 N$19607 N$19828 N$19830 "Waveguide Crossing" sch_x=-238 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5095 N$19609 N$19611 N$19832 N$19834 "Waveguide Crossing" sch_x=-238 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5096 N$19613 N$19615 N$19836 N$19838 "Waveguide Crossing" sch_x=-238 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5097 N$19617 N$19619 N$19840 N$19842 "Waveguide Crossing" sch_x=-238 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5098 N$19621 N$19623 N$19844 N$19846 "Waveguide Crossing" sch_x=-238 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5099 N$19625 N$19627 N$19848 N$19850 "Waveguide Crossing" sch_x=-238 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5100 N$19629 N$19631 N$19852 N$19854 "Waveguide Crossing" sch_x=-238 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5101 N$19633 N$19635 N$19856 N$19858 "Waveguide Crossing" sch_x=-238 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5102 N$19637 N$19639 N$19860 N$19862 "Waveguide Crossing" sch_x=-238 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5103 N$19641 N$19643 N$19864 N$19866 "Waveguide Crossing" sch_x=-238 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5104 N$19645 N$19647 N$19868 N$19870 "Waveguide Crossing" sch_x=-238 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5105 N$19649 N$19651 N$19872 N$19874 "Waveguide Crossing" sch_x=-238 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5106 N$19653 N$19655 N$19876 N$19878 "Waveguide Crossing" sch_x=-238 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5107 N$19657 N$19659 N$19880 N$19882 "Waveguide Crossing" sch_x=-238 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5108 N$19661 N$19663 N$19884 N$19886 "Waveguide Crossing" sch_x=-238 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5109 N$19665 N$19667 N$19888 N$19890 "Waveguide Crossing" sch_x=-238 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5110 N$19669 N$19671 N$19892 N$19894 "Waveguide Crossing" sch_x=-238 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5111 N$19673 N$19675 N$19896 N$19898 "Waveguide Crossing" sch_x=-238 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5112 N$19677 N$19679 N$19900 N$19902 "Waveguide Crossing" sch_x=-238 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5113 N$19681 N$19683 N$19904 N$19906 "Waveguide Crossing" sch_x=-238 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5114 N$19685 N$19687 N$19908 N$19910 "Waveguide Crossing" sch_x=-238 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5115 N$19689 N$19691 N$19912 N$19914 "Waveguide Crossing" sch_x=-238 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5116 N$19693 N$19695 N$19916 N$19918 "Waveguide Crossing" sch_x=-238 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5117 N$19697 N$19699 N$19920 N$19922 "Waveguide Crossing" sch_x=-238 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5118 N$19701 N$19703 N$19924 N$19926 "Waveguide Crossing" sch_x=-238 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5119 N$19705 N$19707 N$19928 N$19930 "Waveguide Crossing" sch_x=-238 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5120 N$19709 N$19711 N$19932 N$19934 "Waveguide Crossing" sch_x=-238 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5121 N$19713 N$19715 N$19936 N$19938 "Waveguide Crossing" sch_x=-238 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5122 N$19717 N$19719 N$19940 N$19942 "Waveguide Crossing" sch_x=-238 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5123 N$19721 N$19723 N$19944 N$19946 "Waveguide Crossing" sch_x=-238 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5124 N$19725 N$19727 N$19948 N$19950 "Waveguide Crossing" sch_x=-238 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5125 N$19729 N$19731 N$19952 N$19954 "Waveguide Crossing" sch_x=-238 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5126 N$19733 N$19735 N$19956 N$19958 "Waveguide Crossing" sch_x=-238 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5127 N$19737 N$19739 N$19960 N$19962 "Waveguide Crossing" sch_x=-238 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5128 N$19741 N$19743 N$19964 N$19966 "Waveguide Crossing" sch_x=-238 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5129 N$19745 N$19747 N$19968 N$19970 "Waveguide Crossing" sch_x=-238 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5130 N$19749 N$19751 N$19972 N$19974 "Waveguide Crossing" sch_x=-238 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5131 N$19753 N$19755 N$19976 N$19978 "Waveguide Crossing" sch_x=-238 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5132 N$19757 N$19759 N$19980 N$19982 "Waveguide Crossing" sch_x=-238 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5133 N$19761 N$19763 N$19984 N$19986 "Waveguide Crossing" sch_x=-238 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5134 N$19765 N$19767 N$19988 N$19990 "Waveguide Crossing" sch_x=-238 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5135 N$19769 N$19771 N$19992 N$19994 "Waveguide Crossing" sch_x=-238 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5136 N$19773 N$19775 N$19996 N$19998 "Waveguide Crossing" sch_x=-238 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5137 N$19777 N$19779 N$20000 N$20002 "Waveguide Crossing" sch_x=-238 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5138 N$19781 N$19783 N$20004 N$20006 "Waveguide Crossing" sch_x=-238 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5139 N$19785 N$19787 N$20008 N$20010 "Waveguide Crossing" sch_x=-238 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5140 N$19789 N$19791 N$20012 N$20014 "Waveguide Crossing" sch_x=-238 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5141 N$19793 N$19795 N$20016 N$20018 "Waveguide Crossing" sch_x=-238 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5142 N$19797 N$19799 N$20020 N$20022 "Waveguide Crossing" sch_x=-238 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5143 N$19801 N$19803 N$20024 N$20026 "Waveguide Crossing" sch_x=-238 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5144 N$19805 N$19807 N$20028 N$20030 "Waveguide Crossing" sch_x=-238 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5145 N$19809 N$19811 N$20032 N$20034 "Waveguide Crossing" sch_x=-238 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5146 N$19813 N$19815 N$20036 N$20038 "Waveguide Crossing" sch_x=-238 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5147 N$19817 N$19819 N$20040 N$20042 "Waveguide Crossing" sch_x=-238 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5148 N$19821 N$19823 N$20044 N$26221 "Waveguide Crossing" sch_x=-238 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5149 N$19825 N$19827 N$26001 N$20046 "Waveguide Crossing" sch_x=-236 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5150 N$19829 N$19831 N$20048 N$20050 "Waveguide Crossing" sch_x=-236 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5151 N$19833 N$19835 N$20052 N$20054 "Waveguide Crossing" sch_x=-236 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5152 N$19837 N$19839 N$20056 N$20058 "Waveguide Crossing" sch_x=-236 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5153 N$19841 N$19843 N$20060 N$20062 "Waveguide Crossing" sch_x=-236 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5154 N$19845 N$19847 N$20064 N$20066 "Waveguide Crossing" sch_x=-236 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5155 N$19849 N$19851 N$20068 N$20070 "Waveguide Crossing" sch_x=-236 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5156 N$19853 N$19855 N$20072 N$20074 "Waveguide Crossing" sch_x=-236 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5157 N$19857 N$19859 N$20076 N$20078 "Waveguide Crossing" sch_x=-236 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5158 N$19861 N$19863 N$20080 N$20082 "Waveguide Crossing" sch_x=-236 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5159 N$19865 N$19867 N$20084 N$20086 "Waveguide Crossing" sch_x=-236 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5160 N$19869 N$19871 N$20088 N$20090 "Waveguide Crossing" sch_x=-236 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5161 N$19873 N$19875 N$20092 N$20094 "Waveguide Crossing" sch_x=-236 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5162 N$19877 N$19879 N$20096 N$20098 "Waveguide Crossing" sch_x=-236 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5163 N$19881 N$19883 N$20100 N$20102 "Waveguide Crossing" sch_x=-236 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5164 N$19885 N$19887 N$20104 N$20106 "Waveguide Crossing" sch_x=-236 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5165 N$19889 N$19891 N$20108 N$20110 "Waveguide Crossing" sch_x=-236 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5166 N$19893 N$19895 N$20112 N$20114 "Waveguide Crossing" sch_x=-236 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5167 N$19897 N$19899 N$20116 N$20118 "Waveguide Crossing" sch_x=-236 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5168 N$19901 N$19903 N$20120 N$20122 "Waveguide Crossing" sch_x=-236 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5169 N$19905 N$19907 N$20124 N$20126 "Waveguide Crossing" sch_x=-236 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5170 N$19909 N$19911 N$20128 N$20130 "Waveguide Crossing" sch_x=-236 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5171 N$19913 N$19915 N$20132 N$20134 "Waveguide Crossing" sch_x=-236 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5172 N$19917 N$19919 N$20136 N$20138 "Waveguide Crossing" sch_x=-236 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5173 N$19921 N$19923 N$20140 N$20142 "Waveguide Crossing" sch_x=-236 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5174 N$19925 N$19927 N$20144 N$20146 "Waveguide Crossing" sch_x=-236 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5175 N$19929 N$19931 N$20148 N$20150 "Waveguide Crossing" sch_x=-236 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5176 N$19933 N$19935 N$20152 N$20154 "Waveguide Crossing" sch_x=-236 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5177 N$19937 N$19939 N$20156 N$20158 "Waveguide Crossing" sch_x=-236 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5178 N$19941 N$19943 N$20160 N$20162 "Waveguide Crossing" sch_x=-236 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5179 N$19945 N$19947 N$20164 N$20166 "Waveguide Crossing" sch_x=-236 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5180 N$19949 N$19951 N$20168 N$20170 "Waveguide Crossing" sch_x=-236 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5181 N$19953 N$19955 N$20172 N$20174 "Waveguide Crossing" sch_x=-236 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5182 N$19957 N$19959 N$20176 N$20178 "Waveguide Crossing" sch_x=-236 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5183 N$19961 N$19963 N$20180 N$20182 "Waveguide Crossing" sch_x=-236 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5184 N$19965 N$19967 N$20184 N$20186 "Waveguide Crossing" sch_x=-236 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5185 N$19969 N$19971 N$20188 N$20190 "Waveguide Crossing" sch_x=-236 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5186 N$19973 N$19975 N$20192 N$20194 "Waveguide Crossing" sch_x=-236 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5187 N$19977 N$19979 N$20196 N$20198 "Waveguide Crossing" sch_x=-236 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5188 N$19981 N$19983 N$20200 N$20202 "Waveguide Crossing" sch_x=-236 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5189 N$19985 N$19987 N$20204 N$20206 "Waveguide Crossing" sch_x=-236 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5190 N$19989 N$19991 N$20208 N$20210 "Waveguide Crossing" sch_x=-236 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5191 N$19993 N$19995 N$20212 N$20214 "Waveguide Crossing" sch_x=-236 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5192 N$19997 N$19999 N$20216 N$20218 "Waveguide Crossing" sch_x=-236 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5193 N$20001 N$20003 N$20220 N$20222 "Waveguide Crossing" sch_x=-236 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5194 N$20005 N$20007 N$20224 N$20226 "Waveguide Crossing" sch_x=-236 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5195 N$20009 N$20011 N$20228 N$20230 "Waveguide Crossing" sch_x=-236 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5196 N$20013 N$20015 N$20232 N$20234 "Waveguide Crossing" sch_x=-236 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5197 N$20017 N$20019 N$20236 N$20238 "Waveguide Crossing" sch_x=-236 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5198 N$20021 N$20023 N$20240 N$20242 "Waveguide Crossing" sch_x=-236 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5199 N$20025 N$20027 N$20244 N$20246 "Waveguide Crossing" sch_x=-236 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5200 N$20029 N$20031 N$20248 N$20250 "Waveguide Crossing" sch_x=-236 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5201 N$20033 N$20035 N$20252 N$20254 "Waveguide Crossing" sch_x=-236 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5202 N$20037 N$20039 N$20256 N$20258 "Waveguide Crossing" sch_x=-236 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5203 N$20041 N$20043 N$20260 N$26219 "Waveguide Crossing" sch_x=-236 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5204 N$20045 N$20047 N$26003 N$20262 "Waveguide Crossing" sch_x=-234 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5205 N$20049 N$20051 N$20264 N$20266 "Waveguide Crossing" sch_x=-234 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5206 N$20053 N$20055 N$20268 N$20270 "Waveguide Crossing" sch_x=-234 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5207 N$20057 N$20059 N$20272 N$20274 "Waveguide Crossing" sch_x=-234 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5208 N$20061 N$20063 N$20276 N$20278 "Waveguide Crossing" sch_x=-234 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5209 N$20065 N$20067 N$20280 N$20282 "Waveguide Crossing" sch_x=-234 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5210 N$20069 N$20071 N$20284 N$20286 "Waveguide Crossing" sch_x=-234 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5211 N$20073 N$20075 N$20288 N$20290 "Waveguide Crossing" sch_x=-234 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5212 N$20077 N$20079 N$20292 N$20294 "Waveguide Crossing" sch_x=-234 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5213 N$20081 N$20083 N$20296 N$20298 "Waveguide Crossing" sch_x=-234 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5214 N$20085 N$20087 N$20300 N$20302 "Waveguide Crossing" sch_x=-234 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5215 N$20089 N$20091 N$20304 N$20306 "Waveguide Crossing" sch_x=-234 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5216 N$20093 N$20095 N$20308 N$20310 "Waveguide Crossing" sch_x=-234 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5217 N$20097 N$20099 N$20312 N$20314 "Waveguide Crossing" sch_x=-234 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5218 N$20101 N$20103 N$20316 N$20318 "Waveguide Crossing" sch_x=-234 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5219 N$20105 N$20107 N$20320 N$20322 "Waveguide Crossing" sch_x=-234 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5220 N$20109 N$20111 N$20324 N$20326 "Waveguide Crossing" sch_x=-234 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5221 N$20113 N$20115 N$20328 N$20330 "Waveguide Crossing" sch_x=-234 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5222 N$20117 N$20119 N$20332 N$20334 "Waveguide Crossing" sch_x=-234 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5223 N$20121 N$20123 N$20336 N$20338 "Waveguide Crossing" sch_x=-234 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5224 N$20125 N$20127 N$20340 N$20342 "Waveguide Crossing" sch_x=-234 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5225 N$20129 N$20131 N$20344 N$20346 "Waveguide Crossing" sch_x=-234 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5226 N$20133 N$20135 N$20348 N$20350 "Waveguide Crossing" sch_x=-234 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5227 N$20137 N$20139 N$20352 N$20354 "Waveguide Crossing" sch_x=-234 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5228 N$20141 N$20143 N$20356 N$20358 "Waveguide Crossing" sch_x=-234 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5229 N$20145 N$20147 N$20360 N$20362 "Waveguide Crossing" sch_x=-234 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5230 N$20149 N$20151 N$20364 N$20366 "Waveguide Crossing" sch_x=-234 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5231 N$20153 N$20155 N$20368 N$20370 "Waveguide Crossing" sch_x=-234 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5232 N$20157 N$20159 N$20372 N$20374 "Waveguide Crossing" sch_x=-234 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5233 N$20161 N$20163 N$20376 N$20378 "Waveguide Crossing" sch_x=-234 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5234 N$20165 N$20167 N$20380 N$20382 "Waveguide Crossing" sch_x=-234 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5235 N$20169 N$20171 N$20384 N$20386 "Waveguide Crossing" sch_x=-234 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5236 N$20173 N$20175 N$20388 N$20390 "Waveguide Crossing" sch_x=-234 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5237 N$20177 N$20179 N$20392 N$20394 "Waveguide Crossing" sch_x=-234 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5238 N$20181 N$20183 N$20396 N$20398 "Waveguide Crossing" sch_x=-234 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5239 N$20185 N$20187 N$20400 N$20402 "Waveguide Crossing" sch_x=-234 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5240 N$20189 N$20191 N$20404 N$20406 "Waveguide Crossing" sch_x=-234 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5241 N$20193 N$20195 N$20408 N$20410 "Waveguide Crossing" sch_x=-234 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5242 N$20197 N$20199 N$20412 N$20414 "Waveguide Crossing" sch_x=-234 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5243 N$20201 N$20203 N$20416 N$20418 "Waveguide Crossing" sch_x=-234 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5244 N$20205 N$20207 N$20420 N$20422 "Waveguide Crossing" sch_x=-234 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5245 N$20209 N$20211 N$20424 N$20426 "Waveguide Crossing" sch_x=-234 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5246 N$20213 N$20215 N$20428 N$20430 "Waveguide Crossing" sch_x=-234 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5247 N$20217 N$20219 N$20432 N$20434 "Waveguide Crossing" sch_x=-234 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5248 N$20221 N$20223 N$20436 N$20438 "Waveguide Crossing" sch_x=-234 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5249 N$20225 N$20227 N$20440 N$20442 "Waveguide Crossing" sch_x=-234 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5250 N$20229 N$20231 N$20444 N$20446 "Waveguide Crossing" sch_x=-234 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5251 N$20233 N$20235 N$20448 N$20450 "Waveguide Crossing" sch_x=-234 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5252 N$20237 N$20239 N$20452 N$20454 "Waveguide Crossing" sch_x=-234 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5253 N$20241 N$20243 N$20456 N$20458 "Waveguide Crossing" sch_x=-234 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5254 N$20245 N$20247 N$20460 N$20462 "Waveguide Crossing" sch_x=-234 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5255 N$20249 N$20251 N$20464 N$20466 "Waveguide Crossing" sch_x=-234 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5256 N$20253 N$20255 N$20468 N$20470 "Waveguide Crossing" sch_x=-234 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5257 N$20257 N$20259 N$20472 N$26217 "Waveguide Crossing" sch_x=-234 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5258 N$20261 N$20263 N$26005 N$20474 "Waveguide Crossing" sch_x=-232 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5259 N$20265 N$20267 N$20476 N$20478 "Waveguide Crossing" sch_x=-232 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5260 N$20269 N$20271 N$20480 N$20482 "Waveguide Crossing" sch_x=-232 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5261 N$20273 N$20275 N$20484 N$20486 "Waveguide Crossing" sch_x=-232 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5262 N$20277 N$20279 N$20488 N$20490 "Waveguide Crossing" sch_x=-232 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5263 N$20281 N$20283 N$20492 N$20494 "Waveguide Crossing" sch_x=-232 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5264 N$20285 N$20287 N$20496 N$20498 "Waveguide Crossing" sch_x=-232 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5265 N$20289 N$20291 N$20500 N$20502 "Waveguide Crossing" sch_x=-232 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5266 N$20293 N$20295 N$20504 N$20506 "Waveguide Crossing" sch_x=-232 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5267 N$20297 N$20299 N$20508 N$20510 "Waveguide Crossing" sch_x=-232 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5268 N$20301 N$20303 N$20512 N$20514 "Waveguide Crossing" sch_x=-232 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5269 N$20305 N$20307 N$20516 N$20518 "Waveguide Crossing" sch_x=-232 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5270 N$20309 N$20311 N$20520 N$20522 "Waveguide Crossing" sch_x=-232 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5271 N$20313 N$20315 N$20524 N$20526 "Waveguide Crossing" sch_x=-232 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5272 N$20317 N$20319 N$20528 N$20530 "Waveguide Crossing" sch_x=-232 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5273 N$20321 N$20323 N$20532 N$20534 "Waveguide Crossing" sch_x=-232 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5274 N$20325 N$20327 N$20536 N$20538 "Waveguide Crossing" sch_x=-232 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5275 N$20329 N$20331 N$20540 N$20542 "Waveguide Crossing" sch_x=-232 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5276 N$20333 N$20335 N$20544 N$20546 "Waveguide Crossing" sch_x=-232 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5277 N$20337 N$20339 N$20548 N$20550 "Waveguide Crossing" sch_x=-232 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5278 N$20341 N$20343 N$20552 N$20554 "Waveguide Crossing" sch_x=-232 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5279 N$20345 N$20347 N$20556 N$20558 "Waveguide Crossing" sch_x=-232 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5280 N$20349 N$20351 N$20560 N$20562 "Waveguide Crossing" sch_x=-232 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5281 N$20353 N$20355 N$20564 N$20566 "Waveguide Crossing" sch_x=-232 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5282 N$20357 N$20359 N$20568 N$20570 "Waveguide Crossing" sch_x=-232 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5283 N$20361 N$20363 N$20572 N$20574 "Waveguide Crossing" sch_x=-232 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5284 N$20365 N$20367 N$20576 N$20578 "Waveguide Crossing" sch_x=-232 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5285 N$20369 N$20371 N$20580 N$20582 "Waveguide Crossing" sch_x=-232 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5286 N$20373 N$20375 N$20584 N$20586 "Waveguide Crossing" sch_x=-232 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5287 N$20377 N$20379 N$20588 N$20590 "Waveguide Crossing" sch_x=-232 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5288 N$20381 N$20383 N$20592 N$20594 "Waveguide Crossing" sch_x=-232 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5289 N$20385 N$20387 N$20596 N$20598 "Waveguide Crossing" sch_x=-232 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5290 N$20389 N$20391 N$20600 N$20602 "Waveguide Crossing" sch_x=-232 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5291 N$20393 N$20395 N$20604 N$20606 "Waveguide Crossing" sch_x=-232 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5292 N$20397 N$20399 N$20608 N$20610 "Waveguide Crossing" sch_x=-232 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5293 N$20401 N$20403 N$20612 N$20614 "Waveguide Crossing" sch_x=-232 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5294 N$20405 N$20407 N$20616 N$20618 "Waveguide Crossing" sch_x=-232 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5295 N$20409 N$20411 N$20620 N$20622 "Waveguide Crossing" sch_x=-232 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5296 N$20413 N$20415 N$20624 N$20626 "Waveguide Crossing" sch_x=-232 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5297 N$20417 N$20419 N$20628 N$20630 "Waveguide Crossing" sch_x=-232 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5298 N$20421 N$20423 N$20632 N$20634 "Waveguide Crossing" sch_x=-232 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5299 N$20425 N$20427 N$20636 N$20638 "Waveguide Crossing" sch_x=-232 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5300 N$20429 N$20431 N$20640 N$20642 "Waveguide Crossing" sch_x=-232 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5301 N$20433 N$20435 N$20644 N$20646 "Waveguide Crossing" sch_x=-232 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5302 N$20437 N$20439 N$20648 N$20650 "Waveguide Crossing" sch_x=-232 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5303 N$20441 N$20443 N$20652 N$20654 "Waveguide Crossing" sch_x=-232 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5304 N$20445 N$20447 N$20656 N$20658 "Waveguide Crossing" sch_x=-232 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5305 N$20449 N$20451 N$20660 N$20662 "Waveguide Crossing" sch_x=-232 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5306 N$20453 N$20455 N$20664 N$20666 "Waveguide Crossing" sch_x=-232 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5307 N$20457 N$20459 N$20668 N$20670 "Waveguide Crossing" sch_x=-232 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5308 N$20461 N$20463 N$20672 N$20674 "Waveguide Crossing" sch_x=-232 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5309 N$20465 N$20467 N$20676 N$20678 "Waveguide Crossing" sch_x=-232 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5310 N$20469 N$20471 N$20680 N$26215 "Waveguide Crossing" sch_x=-232 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5311 N$20473 N$20475 N$26007 N$20682 "Waveguide Crossing" sch_x=-230 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5312 N$20477 N$20479 N$20684 N$20686 "Waveguide Crossing" sch_x=-230 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5313 N$20481 N$20483 N$20688 N$20690 "Waveguide Crossing" sch_x=-230 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5314 N$20485 N$20487 N$20692 N$20694 "Waveguide Crossing" sch_x=-230 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5315 N$20489 N$20491 N$20696 N$20698 "Waveguide Crossing" sch_x=-230 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5316 N$20493 N$20495 N$20700 N$20702 "Waveguide Crossing" sch_x=-230 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5317 N$20497 N$20499 N$20704 N$20706 "Waveguide Crossing" sch_x=-230 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5318 N$20501 N$20503 N$20708 N$20710 "Waveguide Crossing" sch_x=-230 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5319 N$20505 N$20507 N$20712 N$20714 "Waveguide Crossing" sch_x=-230 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5320 N$20509 N$20511 N$20716 N$20718 "Waveguide Crossing" sch_x=-230 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5321 N$20513 N$20515 N$20720 N$20722 "Waveguide Crossing" sch_x=-230 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5322 N$20517 N$20519 N$20724 N$20726 "Waveguide Crossing" sch_x=-230 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5323 N$20521 N$20523 N$20728 N$20730 "Waveguide Crossing" sch_x=-230 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5324 N$20525 N$20527 N$20732 N$20734 "Waveguide Crossing" sch_x=-230 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5325 N$20529 N$20531 N$20736 N$20738 "Waveguide Crossing" sch_x=-230 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5326 N$20533 N$20535 N$20740 N$20742 "Waveguide Crossing" sch_x=-230 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5327 N$20537 N$20539 N$20744 N$20746 "Waveguide Crossing" sch_x=-230 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5328 N$20541 N$20543 N$20748 N$20750 "Waveguide Crossing" sch_x=-230 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5329 N$20545 N$20547 N$20752 N$20754 "Waveguide Crossing" sch_x=-230 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5330 N$20549 N$20551 N$20756 N$20758 "Waveguide Crossing" sch_x=-230 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5331 N$20553 N$20555 N$20760 N$20762 "Waveguide Crossing" sch_x=-230 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5332 N$20557 N$20559 N$20764 N$20766 "Waveguide Crossing" sch_x=-230 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5333 N$20561 N$20563 N$20768 N$20770 "Waveguide Crossing" sch_x=-230 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5334 N$20565 N$20567 N$20772 N$20774 "Waveguide Crossing" sch_x=-230 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5335 N$20569 N$20571 N$20776 N$20778 "Waveguide Crossing" sch_x=-230 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5336 N$20573 N$20575 N$20780 N$20782 "Waveguide Crossing" sch_x=-230 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5337 N$20577 N$20579 N$20784 N$20786 "Waveguide Crossing" sch_x=-230 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5338 N$20581 N$20583 N$20788 N$20790 "Waveguide Crossing" sch_x=-230 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5339 N$20585 N$20587 N$20792 N$20794 "Waveguide Crossing" sch_x=-230 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5340 N$20589 N$20591 N$20796 N$20798 "Waveguide Crossing" sch_x=-230 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5341 N$20593 N$20595 N$20800 N$20802 "Waveguide Crossing" sch_x=-230 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5342 N$20597 N$20599 N$20804 N$20806 "Waveguide Crossing" sch_x=-230 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5343 N$20601 N$20603 N$20808 N$20810 "Waveguide Crossing" sch_x=-230 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5344 N$20605 N$20607 N$20812 N$20814 "Waveguide Crossing" sch_x=-230 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5345 N$20609 N$20611 N$20816 N$20818 "Waveguide Crossing" sch_x=-230 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5346 N$20613 N$20615 N$20820 N$20822 "Waveguide Crossing" sch_x=-230 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5347 N$20617 N$20619 N$20824 N$20826 "Waveguide Crossing" sch_x=-230 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5348 N$20621 N$20623 N$20828 N$20830 "Waveguide Crossing" sch_x=-230 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5349 N$20625 N$20627 N$20832 N$20834 "Waveguide Crossing" sch_x=-230 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5350 N$20629 N$20631 N$20836 N$20838 "Waveguide Crossing" sch_x=-230 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5351 N$20633 N$20635 N$20840 N$20842 "Waveguide Crossing" sch_x=-230 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5352 N$20637 N$20639 N$20844 N$20846 "Waveguide Crossing" sch_x=-230 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5353 N$20641 N$20643 N$20848 N$20850 "Waveguide Crossing" sch_x=-230 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5354 N$20645 N$20647 N$20852 N$20854 "Waveguide Crossing" sch_x=-230 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5355 N$20649 N$20651 N$20856 N$20858 "Waveguide Crossing" sch_x=-230 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5356 N$20653 N$20655 N$20860 N$20862 "Waveguide Crossing" sch_x=-230 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5357 N$20657 N$20659 N$20864 N$20866 "Waveguide Crossing" sch_x=-230 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5358 N$20661 N$20663 N$20868 N$20870 "Waveguide Crossing" sch_x=-230 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5359 N$20665 N$20667 N$20872 N$20874 "Waveguide Crossing" sch_x=-230 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5360 N$20669 N$20671 N$20876 N$20878 "Waveguide Crossing" sch_x=-230 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5361 N$20673 N$20675 N$20880 N$20882 "Waveguide Crossing" sch_x=-230 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5362 N$20677 N$20679 N$20884 N$26213 "Waveguide Crossing" sch_x=-230 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5363 N$20681 N$20683 N$26009 N$20886 "Waveguide Crossing" sch_x=-228 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5364 N$20685 N$20687 N$20888 N$20890 "Waveguide Crossing" sch_x=-228 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5365 N$20689 N$20691 N$20892 N$20894 "Waveguide Crossing" sch_x=-228 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5366 N$20693 N$20695 N$20896 N$20898 "Waveguide Crossing" sch_x=-228 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5367 N$20697 N$20699 N$20900 N$20902 "Waveguide Crossing" sch_x=-228 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5368 N$20701 N$20703 N$20904 N$20906 "Waveguide Crossing" sch_x=-228 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5369 N$20705 N$20707 N$20908 N$20910 "Waveguide Crossing" sch_x=-228 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5370 N$20709 N$20711 N$20912 N$20914 "Waveguide Crossing" sch_x=-228 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5371 N$20713 N$20715 N$20916 N$20918 "Waveguide Crossing" sch_x=-228 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5372 N$20717 N$20719 N$20920 N$20922 "Waveguide Crossing" sch_x=-228 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5373 N$20721 N$20723 N$20924 N$20926 "Waveguide Crossing" sch_x=-228 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5374 N$20725 N$20727 N$20928 N$20930 "Waveguide Crossing" sch_x=-228 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5375 N$20729 N$20731 N$20932 N$20934 "Waveguide Crossing" sch_x=-228 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5376 N$20733 N$20735 N$20936 N$20938 "Waveguide Crossing" sch_x=-228 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5377 N$20737 N$20739 N$20940 N$20942 "Waveguide Crossing" sch_x=-228 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5378 N$20741 N$20743 N$20944 N$20946 "Waveguide Crossing" sch_x=-228 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5379 N$20745 N$20747 N$20948 N$20950 "Waveguide Crossing" sch_x=-228 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5380 N$20749 N$20751 N$20952 N$20954 "Waveguide Crossing" sch_x=-228 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5381 N$20753 N$20755 N$20956 N$20958 "Waveguide Crossing" sch_x=-228 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5382 N$20757 N$20759 N$20960 N$20962 "Waveguide Crossing" sch_x=-228 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5383 N$20761 N$20763 N$20964 N$20966 "Waveguide Crossing" sch_x=-228 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5384 N$20765 N$20767 N$20968 N$20970 "Waveguide Crossing" sch_x=-228 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5385 N$20769 N$20771 N$20972 N$20974 "Waveguide Crossing" sch_x=-228 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5386 N$20773 N$20775 N$20976 N$20978 "Waveguide Crossing" sch_x=-228 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5387 N$20777 N$20779 N$20980 N$20982 "Waveguide Crossing" sch_x=-228 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5388 N$20781 N$20783 N$20984 N$20986 "Waveguide Crossing" sch_x=-228 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5389 N$20785 N$20787 N$20988 N$20990 "Waveguide Crossing" sch_x=-228 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5390 N$20789 N$20791 N$20992 N$20994 "Waveguide Crossing" sch_x=-228 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5391 N$20793 N$20795 N$20996 N$20998 "Waveguide Crossing" sch_x=-228 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5392 N$20797 N$20799 N$21000 N$21002 "Waveguide Crossing" sch_x=-228 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5393 N$20801 N$20803 N$21004 N$21006 "Waveguide Crossing" sch_x=-228 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5394 N$20805 N$20807 N$21008 N$21010 "Waveguide Crossing" sch_x=-228 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5395 N$20809 N$20811 N$21012 N$21014 "Waveguide Crossing" sch_x=-228 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5396 N$20813 N$20815 N$21016 N$21018 "Waveguide Crossing" sch_x=-228 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5397 N$20817 N$20819 N$21020 N$21022 "Waveguide Crossing" sch_x=-228 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5398 N$20821 N$20823 N$21024 N$21026 "Waveguide Crossing" sch_x=-228 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5399 N$20825 N$20827 N$21028 N$21030 "Waveguide Crossing" sch_x=-228 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5400 N$20829 N$20831 N$21032 N$21034 "Waveguide Crossing" sch_x=-228 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5401 N$20833 N$20835 N$21036 N$21038 "Waveguide Crossing" sch_x=-228 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5402 N$20837 N$20839 N$21040 N$21042 "Waveguide Crossing" sch_x=-228 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5403 N$20841 N$20843 N$21044 N$21046 "Waveguide Crossing" sch_x=-228 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5404 N$20845 N$20847 N$21048 N$21050 "Waveguide Crossing" sch_x=-228 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5405 N$20849 N$20851 N$21052 N$21054 "Waveguide Crossing" sch_x=-228 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5406 N$20853 N$20855 N$21056 N$21058 "Waveguide Crossing" sch_x=-228 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5407 N$20857 N$20859 N$21060 N$21062 "Waveguide Crossing" sch_x=-228 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5408 N$20861 N$20863 N$21064 N$21066 "Waveguide Crossing" sch_x=-228 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5409 N$20865 N$20867 N$21068 N$21070 "Waveguide Crossing" sch_x=-228 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5410 N$20869 N$20871 N$21072 N$21074 "Waveguide Crossing" sch_x=-228 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5411 N$20873 N$20875 N$21076 N$21078 "Waveguide Crossing" sch_x=-228 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5412 N$20877 N$20879 N$21080 N$21082 "Waveguide Crossing" sch_x=-228 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5413 N$20881 N$20883 N$21084 N$26211 "Waveguide Crossing" sch_x=-228 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5414 N$20885 N$20887 N$26011 N$21086 "Waveguide Crossing" sch_x=-226 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5415 N$20889 N$20891 N$21088 N$21090 "Waveguide Crossing" sch_x=-226 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5416 N$20893 N$20895 N$21092 N$21094 "Waveguide Crossing" sch_x=-226 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5417 N$20897 N$20899 N$21096 N$21098 "Waveguide Crossing" sch_x=-226 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5418 N$20901 N$20903 N$21100 N$21102 "Waveguide Crossing" sch_x=-226 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5419 N$20905 N$20907 N$21104 N$21106 "Waveguide Crossing" sch_x=-226 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5420 N$20909 N$20911 N$21108 N$21110 "Waveguide Crossing" sch_x=-226 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5421 N$20913 N$20915 N$21112 N$21114 "Waveguide Crossing" sch_x=-226 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5422 N$20917 N$20919 N$21116 N$21118 "Waveguide Crossing" sch_x=-226 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5423 N$20921 N$20923 N$21120 N$21122 "Waveguide Crossing" sch_x=-226 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5424 N$20925 N$20927 N$21124 N$21126 "Waveguide Crossing" sch_x=-226 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5425 N$20929 N$20931 N$21128 N$21130 "Waveguide Crossing" sch_x=-226 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5426 N$20933 N$20935 N$21132 N$21134 "Waveguide Crossing" sch_x=-226 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5427 N$20937 N$20939 N$21136 N$21138 "Waveguide Crossing" sch_x=-226 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5428 N$20941 N$20943 N$21140 N$21142 "Waveguide Crossing" sch_x=-226 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5429 N$20945 N$20947 N$21144 N$21146 "Waveguide Crossing" sch_x=-226 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5430 N$20949 N$20951 N$21148 N$21150 "Waveguide Crossing" sch_x=-226 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5431 N$20953 N$20955 N$21152 N$21154 "Waveguide Crossing" sch_x=-226 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5432 N$20957 N$20959 N$21156 N$21158 "Waveguide Crossing" sch_x=-226 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5433 N$20961 N$20963 N$21160 N$21162 "Waveguide Crossing" sch_x=-226 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5434 N$20965 N$20967 N$21164 N$21166 "Waveguide Crossing" sch_x=-226 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5435 N$20969 N$20971 N$21168 N$21170 "Waveguide Crossing" sch_x=-226 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5436 N$20973 N$20975 N$21172 N$21174 "Waveguide Crossing" sch_x=-226 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5437 N$20977 N$20979 N$21176 N$21178 "Waveguide Crossing" sch_x=-226 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5438 N$20981 N$20983 N$21180 N$21182 "Waveguide Crossing" sch_x=-226 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5439 N$20985 N$20987 N$21184 N$21186 "Waveguide Crossing" sch_x=-226 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5440 N$20989 N$20991 N$21188 N$21190 "Waveguide Crossing" sch_x=-226 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5441 N$20993 N$20995 N$21192 N$21194 "Waveguide Crossing" sch_x=-226 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5442 N$20997 N$20999 N$21196 N$21198 "Waveguide Crossing" sch_x=-226 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5443 N$21001 N$21003 N$21200 N$21202 "Waveguide Crossing" sch_x=-226 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5444 N$21005 N$21007 N$21204 N$21206 "Waveguide Crossing" sch_x=-226 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5445 N$21009 N$21011 N$21208 N$21210 "Waveguide Crossing" sch_x=-226 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5446 N$21013 N$21015 N$21212 N$21214 "Waveguide Crossing" sch_x=-226 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5447 N$21017 N$21019 N$21216 N$21218 "Waveguide Crossing" sch_x=-226 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5448 N$21021 N$21023 N$21220 N$21222 "Waveguide Crossing" sch_x=-226 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5449 N$21025 N$21027 N$21224 N$21226 "Waveguide Crossing" sch_x=-226 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5450 N$21029 N$21031 N$21228 N$21230 "Waveguide Crossing" sch_x=-226 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5451 N$21033 N$21035 N$21232 N$21234 "Waveguide Crossing" sch_x=-226 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5452 N$21037 N$21039 N$21236 N$21238 "Waveguide Crossing" sch_x=-226 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5453 N$21041 N$21043 N$21240 N$21242 "Waveguide Crossing" sch_x=-226 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5454 N$21045 N$21047 N$21244 N$21246 "Waveguide Crossing" sch_x=-226 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5455 N$21049 N$21051 N$21248 N$21250 "Waveguide Crossing" sch_x=-226 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5456 N$21053 N$21055 N$21252 N$21254 "Waveguide Crossing" sch_x=-226 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5457 N$21057 N$21059 N$21256 N$21258 "Waveguide Crossing" sch_x=-226 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5458 N$21061 N$21063 N$21260 N$21262 "Waveguide Crossing" sch_x=-226 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5459 N$21065 N$21067 N$21264 N$21266 "Waveguide Crossing" sch_x=-226 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5460 N$21069 N$21071 N$21268 N$21270 "Waveguide Crossing" sch_x=-226 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5461 N$21073 N$21075 N$21272 N$21274 "Waveguide Crossing" sch_x=-226 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5462 N$21077 N$21079 N$21276 N$21278 "Waveguide Crossing" sch_x=-226 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5463 N$21081 N$21083 N$21280 N$26209 "Waveguide Crossing" sch_x=-226 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5464 N$21085 N$21087 N$26013 N$21282 "Waveguide Crossing" sch_x=-224 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5465 N$21089 N$21091 N$21284 N$21286 "Waveguide Crossing" sch_x=-224 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5466 N$21093 N$21095 N$21288 N$21290 "Waveguide Crossing" sch_x=-224 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5467 N$21097 N$21099 N$21292 N$21294 "Waveguide Crossing" sch_x=-224 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5468 N$21101 N$21103 N$21296 N$21298 "Waveguide Crossing" sch_x=-224 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5469 N$21105 N$21107 N$21300 N$21302 "Waveguide Crossing" sch_x=-224 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5470 N$21109 N$21111 N$21304 N$21306 "Waveguide Crossing" sch_x=-224 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5471 N$21113 N$21115 N$21308 N$21310 "Waveguide Crossing" sch_x=-224 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5472 N$21117 N$21119 N$21312 N$21314 "Waveguide Crossing" sch_x=-224 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5473 N$21121 N$21123 N$21316 N$21318 "Waveguide Crossing" sch_x=-224 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5474 N$21125 N$21127 N$21320 N$21322 "Waveguide Crossing" sch_x=-224 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5475 N$21129 N$21131 N$21324 N$21326 "Waveguide Crossing" sch_x=-224 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5476 N$21133 N$21135 N$21328 N$21330 "Waveguide Crossing" sch_x=-224 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5477 N$21137 N$21139 N$21332 N$21334 "Waveguide Crossing" sch_x=-224 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5478 N$21141 N$21143 N$21336 N$21338 "Waveguide Crossing" sch_x=-224 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5479 N$21145 N$21147 N$21340 N$21342 "Waveguide Crossing" sch_x=-224 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5480 N$21149 N$21151 N$21344 N$21346 "Waveguide Crossing" sch_x=-224 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5481 N$21153 N$21155 N$21348 N$21350 "Waveguide Crossing" sch_x=-224 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5482 N$21157 N$21159 N$21352 N$21354 "Waveguide Crossing" sch_x=-224 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5483 N$21161 N$21163 N$21356 N$21358 "Waveguide Crossing" sch_x=-224 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5484 N$21165 N$21167 N$21360 N$21362 "Waveguide Crossing" sch_x=-224 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5485 N$21169 N$21171 N$21364 N$21366 "Waveguide Crossing" sch_x=-224 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5486 N$21173 N$21175 N$21368 N$21370 "Waveguide Crossing" sch_x=-224 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5487 N$21177 N$21179 N$21372 N$21374 "Waveguide Crossing" sch_x=-224 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5488 N$21181 N$21183 N$21376 N$21378 "Waveguide Crossing" sch_x=-224 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5489 N$21185 N$21187 N$21380 N$21382 "Waveguide Crossing" sch_x=-224 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5490 N$21189 N$21191 N$21384 N$21386 "Waveguide Crossing" sch_x=-224 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5491 N$21193 N$21195 N$21388 N$21390 "Waveguide Crossing" sch_x=-224 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5492 N$21197 N$21199 N$21392 N$21394 "Waveguide Crossing" sch_x=-224 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5493 N$21201 N$21203 N$21396 N$21398 "Waveguide Crossing" sch_x=-224 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5494 N$21205 N$21207 N$21400 N$21402 "Waveguide Crossing" sch_x=-224 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5495 N$21209 N$21211 N$21404 N$21406 "Waveguide Crossing" sch_x=-224 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5496 N$21213 N$21215 N$21408 N$21410 "Waveguide Crossing" sch_x=-224 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5497 N$21217 N$21219 N$21412 N$21414 "Waveguide Crossing" sch_x=-224 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5498 N$21221 N$21223 N$21416 N$21418 "Waveguide Crossing" sch_x=-224 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5499 N$21225 N$21227 N$21420 N$21422 "Waveguide Crossing" sch_x=-224 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5500 N$21229 N$21231 N$21424 N$21426 "Waveguide Crossing" sch_x=-224 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5501 N$21233 N$21235 N$21428 N$21430 "Waveguide Crossing" sch_x=-224 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5502 N$21237 N$21239 N$21432 N$21434 "Waveguide Crossing" sch_x=-224 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5503 N$21241 N$21243 N$21436 N$21438 "Waveguide Crossing" sch_x=-224 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5504 N$21245 N$21247 N$21440 N$21442 "Waveguide Crossing" sch_x=-224 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5505 N$21249 N$21251 N$21444 N$21446 "Waveguide Crossing" sch_x=-224 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5506 N$21253 N$21255 N$21448 N$21450 "Waveguide Crossing" sch_x=-224 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5507 N$21257 N$21259 N$21452 N$21454 "Waveguide Crossing" sch_x=-224 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5508 N$21261 N$21263 N$21456 N$21458 "Waveguide Crossing" sch_x=-224 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5509 N$21265 N$21267 N$21460 N$21462 "Waveguide Crossing" sch_x=-224 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5510 N$21269 N$21271 N$21464 N$21466 "Waveguide Crossing" sch_x=-224 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5511 N$21273 N$21275 N$21468 N$21470 "Waveguide Crossing" sch_x=-224 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5512 N$21277 N$21279 N$21472 N$26207 "Waveguide Crossing" sch_x=-224 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5513 N$21281 N$21283 N$26015 N$21474 "Waveguide Crossing" sch_x=-222 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5514 N$21285 N$21287 N$21476 N$21478 "Waveguide Crossing" sch_x=-222 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5515 N$21289 N$21291 N$21480 N$21482 "Waveguide Crossing" sch_x=-222 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5516 N$21293 N$21295 N$21484 N$21486 "Waveguide Crossing" sch_x=-222 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5517 N$21297 N$21299 N$21488 N$21490 "Waveguide Crossing" sch_x=-222 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5518 N$21301 N$21303 N$21492 N$21494 "Waveguide Crossing" sch_x=-222 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5519 N$21305 N$21307 N$21496 N$21498 "Waveguide Crossing" sch_x=-222 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5520 N$21309 N$21311 N$21500 N$21502 "Waveguide Crossing" sch_x=-222 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5521 N$21313 N$21315 N$21504 N$21506 "Waveguide Crossing" sch_x=-222 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5522 N$21317 N$21319 N$21508 N$21510 "Waveguide Crossing" sch_x=-222 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5523 N$21321 N$21323 N$21512 N$21514 "Waveguide Crossing" sch_x=-222 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5524 N$21325 N$21327 N$21516 N$21518 "Waveguide Crossing" sch_x=-222 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5525 N$21329 N$21331 N$21520 N$21522 "Waveguide Crossing" sch_x=-222 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5526 N$21333 N$21335 N$21524 N$21526 "Waveguide Crossing" sch_x=-222 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5527 N$21337 N$21339 N$21528 N$21530 "Waveguide Crossing" sch_x=-222 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5528 N$21341 N$21343 N$21532 N$21534 "Waveguide Crossing" sch_x=-222 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5529 N$21345 N$21347 N$21536 N$21538 "Waveguide Crossing" sch_x=-222 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5530 N$21349 N$21351 N$21540 N$21542 "Waveguide Crossing" sch_x=-222 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5531 N$21353 N$21355 N$21544 N$21546 "Waveguide Crossing" sch_x=-222 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5532 N$21357 N$21359 N$21548 N$21550 "Waveguide Crossing" sch_x=-222 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5533 N$21361 N$21363 N$21552 N$21554 "Waveguide Crossing" sch_x=-222 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5534 N$21365 N$21367 N$21556 N$21558 "Waveguide Crossing" sch_x=-222 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5535 N$21369 N$21371 N$21560 N$21562 "Waveguide Crossing" sch_x=-222 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5536 N$21373 N$21375 N$21564 N$21566 "Waveguide Crossing" sch_x=-222 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5537 N$21377 N$21379 N$21568 N$21570 "Waveguide Crossing" sch_x=-222 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5538 N$21381 N$21383 N$21572 N$21574 "Waveguide Crossing" sch_x=-222 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5539 N$21385 N$21387 N$21576 N$21578 "Waveguide Crossing" sch_x=-222 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5540 N$21389 N$21391 N$21580 N$21582 "Waveguide Crossing" sch_x=-222 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5541 N$21393 N$21395 N$21584 N$21586 "Waveguide Crossing" sch_x=-222 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5542 N$21397 N$21399 N$21588 N$21590 "Waveguide Crossing" sch_x=-222 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5543 N$21401 N$21403 N$21592 N$21594 "Waveguide Crossing" sch_x=-222 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5544 N$21405 N$21407 N$21596 N$21598 "Waveguide Crossing" sch_x=-222 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5545 N$21409 N$21411 N$21600 N$21602 "Waveguide Crossing" sch_x=-222 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5546 N$21413 N$21415 N$21604 N$21606 "Waveguide Crossing" sch_x=-222 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5547 N$21417 N$21419 N$21608 N$21610 "Waveguide Crossing" sch_x=-222 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5548 N$21421 N$21423 N$21612 N$21614 "Waveguide Crossing" sch_x=-222 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5549 N$21425 N$21427 N$21616 N$21618 "Waveguide Crossing" sch_x=-222 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5550 N$21429 N$21431 N$21620 N$21622 "Waveguide Crossing" sch_x=-222 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5551 N$21433 N$21435 N$21624 N$21626 "Waveguide Crossing" sch_x=-222 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5552 N$21437 N$21439 N$21628 N$21630 "Waveguide Crossing" sch_x=-222 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5553 N$21441 N$21443 N$21632 N$21634 "Waveguide Crossing" sch_x=-222 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5554 N$21445 N$21447 N$21636 N$21638 "Waveguide Crossing" sch_x=-222 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5555 N$21449 N$21451 N$21640 N$21642 "Waveguide Crossing" sch_x=-222 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5556 N$21453 N$21455 N$21644 N$21646 "Waveguide Crossing" sch_x=-222 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5557 N$21457 N$21459 N$21648 N$21650 "Waveguide Crossing" sch_x=-222 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5558 N$21461 N$21463 N$21652 N$21654 "Waveguide Crossing" sch_x=-222 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5559 N$21465 N$21467 N$21656 N$21658 "Waveguide Crossing" sch_x=-222 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5560 N$21469 N$21471 N$21660 N$26205 "Waveguide Crossing" sch_x=-222 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5561 N$21473 N$21475 N$26017 N$21662 "Waveguide Crossing" sch_x=-220 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5562 N$21477 N$21479 N$21664 N$21666 "Waveguide Crossing" sch_x=-220 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5563 N$21481 N$21483 N$21668 N$21670 "Waveguide Crossing" sch_x=-220 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5564 N$21485 N$21487 N$21672 N$21674 "Waveguide Crossing" sch_x=-220 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5565 N$21489 N$21491 N$21676 N$21678 "Waveguide Crossing" sch_x=-220 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5566 N$21493 N$21495 N$21680 N$21682 "Waveguide Crossing" sch_x=-220 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5567 N$21497 N$21499 N$21684 N$21686 "Waveguide Crossing" sch_x=-220 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5568 N$21501 N$21503 N$21688 N$21690 "Waveguide Crossing" sch_x=-220 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5569 N$21505 N$21507 N$21692 N$21694 "Waveguide Crossing" sch_x=-220 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5570 N$21509 N$21511 N$21696 N$21698 "Waveguide Crossing" sch_x=-220 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5571 N$21513 N$21515 N$21700 N$21702 "Waveguide Crossing" sch_x=-220 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5572 N$21517 N$21519 N$21704 N$21706 "Waveguide Crossing" sch_x=-220 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5573 N$21521 N$21523 N$21708 N$21710 "Waveguide Crossing" sch_x=-220 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5574 N$21525 N$21527 N$21712 N$21714 "Waveguide Crossing" sch_x=-220 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5575 N$21529 N$21531 N$21716 N$21718 "Waveguide Crossing" sch_x=-220 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5576 N$21533 N$21535 N$21720 N$21722 "Waveguide Crossing" sch_x=-220 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5577 N$21537 N$21539 N$21724 N$21726 "Waveguide Crossing" sch_x=-220 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5578 N$21541 N$21543 N$21728 N$21730 "Waveguide Crossing" sch_x=-220 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5579 N$21545 N$21547 N$21732 N$21734 "Waveguide Crossing" sch_x=-220 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5580 N$21549 N$21551 N$21736 N$21738 "Waveguide Crossing" sch_x=-220 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5581 N$21553 N$21555 N$21740 N$21742 "Waveguide Crossing" sch_x=-220 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5582 N$21557 N$21559 N$21744 N$21746 "Waveguide Crossing" sch_x=-220 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5583 N$21561 N$21563 N$21748 N$21750 "Waveguide Crossing" sch_x=-220 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5584 N$21565 N$21567 N$21752 N$21754 "Waveguide Crossing" sch_x=-220 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5585 N$21569 N$21571 N$21756 N$21758 "Waveguide Crossing" sch_x=-220 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5586 N$21573 N$21575 N$21760 N$21762 "Waveguide Crossing" sch_x=-220 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5587 N$21577 N$21579 N$21764 N$21766 "Waveguide Crossing" sch_x=-220 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5588 N$21581 N$21583 N$21768 N$21770 "Waveguide Crossing" sch_x=-220 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5589 N$21585 N$21587 N$21772 N$21774 "Waveguide Crossing" sch_x=-220 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5590 N$21589 N$21591 N$21776 N$21778 "Waveguide Crossing" sch_x=-220 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5591 N$21593 N$21595 N$21780 N$21782 "Waveguide Crossing" sch_x=-220 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5592 N$21597 N$21599 N$21784 N$21786 "Waveguide Crossing" sch_x=-220 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5593 N$21601 N$21603 N$21788 N$21790 "Waveguide Crossing" sch_x=-220 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5594 N$21605 N$21607 N$21792 N$21794 "Waveguide Crossing" sch_x=-220 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5595 N$21609 N$21611 N$21796 N$21798 "Waveguide Crossing" sch_x=-220 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5596 N$21613 N$21615 N$21800 N$21802 "Waveguide Crossing" sch_x=-220 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5597 N$21617 N$21619 N$21804 N$21806 "Waveguide Crossing" sch_x=-220 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5598 N$21621 N$21623 N$21808 N$21810 "Waveguide Crossing" sch_x=-220 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5599 N$21625 N$21627 N$21812 N$21814 "Waveguide Crossing" sch_x=-220 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5600 N$21629 N$21631 N$21816 N$21818 "Waveguide Crossing" sch_x=-220 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5601 N$21633 N$21635 N$21820 N$21822 "Waveguide Crossing" sch_x=-220 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5602 N$21637 N$21639 N$21824 N$21826 "Waveguide Crossing" sch_x=-220 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5603 N$21641 N$21643 N$21828 N$21830 "Waveguide Crossing" sch_x=-220 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5604 N$21645 N$21647 N$21832 N$21834 "Waveguide Crossing" sch_x=-220 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5605 N$21649 N$21651 N$21836 N$21838 "Waveguide Crossing" sch_x=-220 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5606 N$21653 N$21655 N$21840 N$21842 "Waveguide Crossing" sch_x=-220 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5607 N$21657 N$21659 N$21844 N$26203 "Waveguide Crossing" sch_x=-220 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5608 N$21661 N$21663 N$26019 N$21846 "Waveguide Crossing" sch_x=-218 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5609 N$21665 N$21667 N$21848 N$21850 "Waveguide Crossing" sch_x=-218 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5610 N$21669 N$21671 N$21852 N$21854 "Waveguide Crossing" sch_x=-218 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5611 N$21673 N$21675 N$21856 N$21858 "Waveguide Crossing" sch_x=-218 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5612 N$21677 N$21679 N$21860 N$21862 "Waveguide Crossing" sch_x=-218 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5613 N$21681 N$21683 N$21864 N$21866 "Waveguide Crossing" sch_x=-218 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5614 N$21685 N$21687 N$21868 N$21870 "Waveguide Crossing" sch_x=-218 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5615 N$21689 N$21691 N$21872 N$21874 "Waveguide Crossing" sch_x=-218 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5616 N$21693 N$21695 N$21876 N$21878 "Waveguide Crossing" sch_x=-218 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5617 N$21697 N$21699 N$21880 N$21882 "Waveguide Crossing" sch_x=-218 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5618 N$21701 N$21703 N$21884 N$21886 "Waveguide Crossing" sch_x=-218 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5619 N$21705 N$21707 N$21888 N$21890 "Waveguide Crossing" sch_x=-218 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5620 N$21709 N$21711 N$21892 N$21894 "Waveguide Crossing" sch_x=-218 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5621 N$21713 N$21715 N$21896 N$21898 "Waveguide Crossing" sch_x=-218 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5622 N$21717 N$21719 N$21900 N$21902 "Waveguide Crossing" sch_x=-218 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5623 N$21721 N$21723 N$21904 N$21906 "Waveguide Crossing" sch_x=-218 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5624 N$21725 N$21727 N$21908 N$21910 "Waveguide Crossing" sch_x=-218 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5625 N$21729 N$21731 N$21912 N$21914 "Waveguide Crossing" sch_x=-218 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5626 N$21733 N$21735 N$21916 N$21918 "Waveguide Crossing" sch_x=-218 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5627 N$21737 N$21739 N$21920 N$21922 "Waveguide Crossing" sch_x=-218 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5628 N$21741 N$21743 N$21924 N$21926 "Waveguide Crossing" sch_x=-218 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5629 N$21745 N$21747 N$21928 N$21930 "Waveguide Crossing" sch_x=-218 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5630 N$21749 N$21751 N$21932 N$21934 "Waveguide Crossing" sch_x=-218 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5631 N$21753 N$21755 N$21936 N$21938 "Waveguide Crossing" sch_x=-218 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5632 N$21757 N$21759 N$21940 N$21942 "Waveguide Crossing" sch_x=-218 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5633 N$21761 N$21763 N$21944 N$21946 "Waveguide Crossing" sch_x=-218 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5634 N$21765 N$21767 N$21948 N$21950 "Waveguide Crossing" sch_x=-218 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5635 N$21769 N$21771 N$21952 N$21954 "Waveguide Crossing" sch_x=-218 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5636 N$21773 N$21775 N$21956 N$21958 "Waveguide Crossing" sch_x=-218 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5637 N$21777 N$21779 N$21960 N$21962 "Waveguide Crossing" sch_x=-218 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5638 N$21781 N$21783 N$21964 N$21966 "Waveguide Crossing" sch_x=-218 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5639 N$21785 N$21787 N$21968 N$21970 "Waveguide Crossing" sch_x=-218 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5640 N$21789 N$21791 N$21972 N$21974 "Waveguide Crossing" sch_x=-218 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5641 N$21793 N$21795 N$21976 N$21978 "Waveguide Crossing" sch_x=-218 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5642 N$21797 N$21799 N$21980 N$21982 "Waveguide Crossing" sch_x=-218 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5643 N$21801 N$21803 N$21984 N$21986 "Waveguide Crossing" sch_x=-218 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5644 N$21805 N$21807 N$21988 N$21990 "Waveguide Crossing" sch_x=-218 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5645 N$21809 N$21811 N$21992 N$21994 "Waveguide Crossing" sch_x=-218 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5646 N$21813 N$21815 N$21996 N$21998 "Waveguide Crossing" sch_x=-218 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5647 N$21817 N$21819 N$22000 N$22002 "Waveguide Crossing" sch_x=-218 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5648 N$21821 N$21823 N$22004 N$22006 "Waveguide Crossing" sch_x=-218 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5649 N$21825 N$21827 N$22008 N$22010 "Waveguide Crossing" sch_x=-218 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5650 N$21829 N$21831 N$22012 N$22014 "Waveguide Crossing" sch_x=-218 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5651 N$21833 N$21835 N$22016 N$22018 "Waveguide Crossing" sch_x=-218 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5652 N$21837 N$21839 N$22020 N$22022 "Waveguide Crossing" sch_x=-218 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5653 N$21841 N$21843 N$22024 N$26201 "Waveguide Crossing" sch_x=-218 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5654 N$21845 N$21847 N$26021 N$22026 "Waveguide Crossing" sch_x=-216 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5655 N$21849 N$21851 N$22028 N$22030 "Waveguide Crossing" sch_x=-216 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5656 N$21853 N$21855 N$22032 N$22034 "Waveguide Crossing" sch_x=-216 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5657 N$21857 N$21859 N$22036 N$22038 "Waveguide Crossing" sch_x=-216 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5658 N$21861 N$21863 N$22040 N$22042 "Waveguide Crossing" sch_x=-216 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5659 N$21865 N$21867 N$22044 N$22046 "Waveguide Crossing" sch_x=-216 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5660 N$21869 N$21871 N$22048 N$22050 "Waveguide Crossing" sch_x=-216 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5661 N$21873 N$21875 N$22052 N$22054 "Waveguide Crossing" sch_x=-216 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5662 N$21877 N$21879 N$22056 N$22058 "Waveguide Crossing" sch_x=-216 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5663 N$21881 N$21883 N$22060 N$22062 "Waveguide Crossing" sch_x=-216 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5664 N$21885 N$21887 N$22064 N$22066 "Waveguide Crossing" sch_x=-216 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5665 N$21889 N$21891 N$22068 N$22070 "Waveguide Crossing" sch_x=-216 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5666 N$21893 N$21895 N$22072 N$22074 "Waveguide Crossing" sch_x=-216 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5667 N$21897 N$21899 N$22076 N$22078 "Waveguide Crossing" sch_x=-216 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5668 N$21901 N$21903 N$22080 N$22082 "Waveguide Crossing" sch_x=-216 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5669 N$21905 N$21907 N$22084 N$22086 "Waveguide Crossing" sch_x=-216 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5670 N$21909 N$21911 N$22088 N$22090 "Waveguide Crossing" sch_x=-216 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5671 N$21913 N$21915 N$22092 N$22094 "Waveguide Crossing" sch_x=-216 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5672 N$21917 N$21919 N$22096 N$22098 "Waveguide Crossing" sch_x=-216 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5673 N$21921 N$21923 N$22100 N$22102 "Waveguide Crossing" sch_x=-216 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5674 N$21925 N$21927 N$22104 N$22106 "Waveguide Crossing" sch_x=-216 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5675 N$21929 N$21931 N$22108 N$22110 "Waveguide Crossing" sch_x=-216 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5676 N$21933 N$21935 N$22112 N$22114 "Waveguide Crossing" sch_x=-216 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5677 N$21937 N$21939 N$22116 N$22118 "Waveguide Crossing" sch_x=-216 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5678 N$21941 N$21943 N$22120 N$22122 "Waveguide Crossing" sch_x=-216 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5679 N$21945 N$21947 N$22124 N$22126 "Waveguide Crossing" sch_x=-216 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5680 N$21949 N$21951 N$22128 N$22130 "Waveguide Crossing" sch_x=-216 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5681 N$21953 N$21955 N$22132 N$22134 "Waveguide Crossing" sch_x=-216 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5682 N$21957 N$21959 N$22136 N$22138 "Waveguide Crossing" sch_x=-216 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5683 N$21961 N$21963 N$22140 N$22142 "Waveguide Crossing" sch_x=-216 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5684 N$21965 N$21967 N$22144 N$22146 "Waveguide Crossing" sch_x=-216 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5685 N$21969 N$21971 N$22148 N$22150 "Waveguide Crossing" sch_x=-216 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5686 N$21973 N$21975 N$22152 N$22154 "Waveguide Crossing" sch_x=-216 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5687 N$21977 N$21979 N$22156 N$22158 "Waveguide Crossing" sch_x=-216 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5688 N$21981 N$21983 N$22160 N$22162 "Waveguide Crossing" sch_x=-216 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5689 N$21985 N$21987 N$22164 N$22166 "Waveguide Crossing" sch_x=-216 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5690 N$21989 N$21991 N$22168 N$22170 "Waveguide Crossing" sch_x=-216 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5691 N$21993 N$21995 N$22172 N$22174 "Waveguide Crossing" sch_x=-216 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5692 N$21997 N$21999 N$22176 N$22178 "Waveguide Crossing" sch_x=-216 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5693 N$22001 N$22003 N$22180 N$22182 "Waveguide Crossing" sch_x=-216 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5694 N$22005 N$22007 N$22184 N$22186 "Waveguide Crossing" sch_x=-216 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5695 N$22009 N$22011 N$22188 N$22190 "Waveguide Crossing" sch_x=-216 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5696 N$22013 N$22015 N$22192 N$22194 "Waveguide Crossing" sch_x=-216 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5697 N$22017 N$22019 N$22196 N$22198 "Waveguide Crossing" sch_x=-216 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5698 N$22021 N$22023 N$22200 N$26199 "Waveguide Crossing" sch_x=-216 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5699 N$22025 N$22027 N$26023 N$22202 "Waveguide Crossing" sch_x=-214 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5700 N$22029 N$22031 N$22204 N$22206 "Waveguide Crossing" sch_x=-214 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5701 N$22033 N$22035 N$22208 N$22210 "Waveguide Crossing" sch_x=-214 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5702 N$22037 N$22039 N$22212 N$22214 "Waveguide Crossing" sch_x=-214 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5703 N$22041 N$22043 N$22216 N$22218 "Waveguide Crossing" sch_x=-214 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5704 N$22045 N$22047 N$22220 N$22222 "Waveguide Crossing" sch_x=-214 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5705 N$22049 N$22051 N$22224 N$22226 "Waveguide Crossing" sch_x=-214 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5706 N$22053 N$22055 N$22228 N$22230 "Waveguide Crossing" sch_x=-214 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5707 N$22057 N$22059 N$22232 N$22234 "Waveguide Crossing" sch_x=-214 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5708 N$22061 N$22063 N$22236 N$22238 "Waveguide Crossing" sch_x=-214 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5709 N$22065 N$22067 N$22240 N$22242 "Waveguide Crossing" sch_x=-214 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5710 N$22069 N$22071 N$22244 N$22246 "Waveguide Crossing" sch_x=-214 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5711 N$22073 N$22075 N$22248 N$22250 "Waveguide Crossing" sch_x=-214 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5712 N$22077 N$22079 N$22252 N$22254 "Waveguide Crossing" sch_x=-214 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5713 N$22081 N$22083 N$22256 N$22258 "Waveguide Crossing" sch_x=-214 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5714 N$22085 N$22087 N$22260 N$22262 "Waveguide Crossing" sch_x=-214 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5715 N$22089 N$22091 N$22264 N$22266 "Waveguide Crossing" sch_x=-214 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5716 N$22093 N$22095 N$22268 N$22270 "Waveguide Crossing" sch_x=-214 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5717 N$22097 N$22099 N$22272 N$22274 "Waveguide Crossing" sch_x=-214 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5718 N$22101 N$22103 N$22276 N$22278 "Waveguide Crossing" sch_x=-214 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5719 N$22105 N$22107 N$22280 N$22282 "Waveguide Crossing" sch_x=-214 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5720 N$22109 N$22111 N$22284 N$22286 "Waveguide Crossing" sch_x=-214 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5721 N$22113 N$22115 N$22288 N$22290 "Waveguide Crossing" sch_x=-214 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5722 N$22117 N$22119 N$22292 N$22294 "Waveguide Crossing" sch_x=-214 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5723 N$22121 N$22123 N$22296 N$22298 "Waveguide Crossing" sch_x=-214 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5724 N$22125 N$22127 N$22300 N$22302 "Waveguide Crossing" sch_x=-214 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5725 N$22129 N$22131 N$22304 N$22306 "Waveguide Crossing" sch_x=-214 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5726 N$22133 N$22135 N$22308 N$22310 "Waveguide Crossing" sch_x=-214 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5727 N$22137 N$22139 N$22312 N$22314 "Waveguide Crossing" sch_x=-214 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5728 N$22141 N$22143 N$22316 N$22318 "Waveguide Crossing" sch_x=-214 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5729 N$22145 N$22147 N$22320 N$22322 "Waveguide Crossing" sch_x=-214 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5730 N$22149 N$22151 N$22324 N$22326 "Waveguide Crossing" sch_x=-214 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5731 N$22153 N$22155 N$22328 N$22330 "Waveguide Crossing" sch_x=-214 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5732 N$22157 N$22159 N$22332 N$22334 "Waveguide Crossing" sch_x=-214 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5733 N$22161 N$22163 N$22336 N$22338 "Waveguide Crossing" sch_x=-214 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5734 N$22165 N$22167 N$22340 N$22342 "Waveguide Crossing" sch_x=-214 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5735 N$22169 N$22171 N$22344 N$22346 "Waveguide Crossing" sch_x=-214 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5736 N$22173 N$22175 N$22348 N$22350 "Waveguide Crossing" sch_x=-214 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5737 N$22177 N$22179 N$22352 N$22354 "Waveguide Crossing" sch_x=-214 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5738 N$22181 N$22183 N$22356 N$22358 "Waveguide Crossing" sch_x=-214 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5739 N$22185 N$22187 N$22360 N$22362 "Waveguide Crossing" sch_x=-214 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5740 N$22189 N$22191 N$22364 N$22366 "Waveguide Crossing" sch_x=-214 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5741 N$22193 N$22195 N$22368 N$22370 "Waveguide Crossing" sch_x=-214 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5742 N$22197 N$22199 N$22372 N$26197 "Waveguide Crossing" sch_x=-214 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5743 N$22201 N$22203 N$26025 N$22374 "Waveguide Crossing" sch_x=-212 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5744 N$22205 N$22207 N$22376 N$22378 "Waveguide Crossing" sch_x=-212 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5745 N$22209 N$22211 N$22380 N$22382 "Waveguide Crossing" sch_x=-212 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5746 N$22213 N$22215 N$22384 N$22386 "Waveguide Crossing" sch_x=-212 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5747 N$22217 N$22219 N$22388 N$22390 "Waveguide Crossing" sch_x=-212 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5748 N$22221 N$22223 N$22392 N$22394 "Waveguide Crossing" sch_x=-212 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5749 N$22225 N$22227 N$22396 N$22398 "Waveguide Crossing" sch_x=-212 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5750 N$22229 N$22231 N$22400 N$22402 "Waveguide Crossing" sch_x=-212 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5751 N$22233 N$22235 N$22404 N$22406 "Waveguide Crossing" sch_x=-212 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5752 N$22237 N$22239 N$22408 N$22410 "Waveguide Crossing" sch_x=-212 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5753 N$22241 N$22243 N$22412 N$22414 "Waveguide Crossing" sch_x=-212 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5754 N$22245 N$22247 N$22416 N$22418 "Waveguide Crossing" sch_x=-212 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5755 N$22249 N$22251 N$22420 N$22422 "Waveguide Crossing" sch_x=-212 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5756 N$22253 N$22255 N$22424 N$22426 "Waveguide Crossing" sch_x=-212 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5757 N$22257 N$22259 N$22428 N$22430 "Waveguide Crossing" sch_x=-212 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5758 N$22261 N$22263 N$22432 N$22434 "Waveguide Crossing" sch_x=-212 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5759 N$22265 N$22267 N$22436 N$22438 "Waveguide Crossing" sch_x=-212 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5760 N$22269 N$22271 N$22440 N$22442 "Waveguide Crossing" sch_x=-212 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5761 N$22273 N$22275 N$22444 N$22446 "Waveguide Crossing" sch_x=-212 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5762 N$22277 N$22279 N$22448 N$22450 "Waveguide Crossing" sch_x=-212 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5763 N$22281 N$22283 N$22452 N$22454 "Waveguide Crossing" sch_x=-212 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5764 N$22285 N$22287 N$22456 N$22458 "Waveguide Crossing" sch_x=-212 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5765 N$22289 N$22291 N$22460 N$22462 "Waveguide Crossing" sch_x=-212 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5766 N$22293 N$22295 N$22464 N$22466 "Waveguide Crossing" sch_x=-212 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5767 N$22297 N$22299 N$22468 N$22470 "Waveguide Crossing" sch_x=-212 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5768 N$22301 N$22303 N$22472 N$22474 "Waveguide Crossing" sch_x=-212 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5769 N$22305 N$22307 N$22476 N$22478 "Waveguide Crossing" sch_x=-212 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5770 N$22309 N$22311 N$22480 N$22482 "Waveguide Crossing" sch_x=-212 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5771 N$22313 N$22315 N$22484 N$22486 "Waveguide Crossing" sch_x=-212 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5772 N$22317 N$22319 N$22488 N$22490 "Waveguide Crossing" sch_x=-212 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5773 N$22321 N$22323 N$22492 N$22494 "Waveguide Crossing" sch_x=-212 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5774 N$22325 N$22327 N$22496 N$22498 "Waveguide Crossing" sch_x=-212 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5775 N$22329 N$22331 N$22500 N$22502 "Waveguide Crossing" sch_x=-212 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5776 N$22333 N$22335 N$22504 N$22506 "Waveguide Crossing" sch_x=-212 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5777 N$22337 N$22339 N$22508 N$22510 "Waveguide Crossing" sch_x=-212 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5778 N$22341 N$22343 N$22512 N$22514 "Waveguide Crossing" sch_x=-212 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5779 N$22345 N$22347 N$22516 N$22518 "Waveguide Crossing" sch_x=-212 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5780 N$22349 N$22351 N$22520 N$22522 "Waveguide Crossing" sch_x=-212 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5781 N$22353 N$22355 N$22524 N$22526 "Waveguide Crossing" sch_x=-212 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5782 N$22357 N$22359 N$22528 N$22530 "Waveguide Crossing" sch_x=-212 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5783 N$22361 N$22363 N$22532 N$22534 "Waveguide Crossing" sch_x=-212 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5784 N$22365 N$22367 N$22536 N$22538 "Waveguide Crossing" sch_x=-212 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5785 N$22369 N$22371 N$22540 N$26195 "Waveguide Crossing" sch_x=-212 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5786 N$22373 N$22375 N$26027 N$22542 "Waveguide Crossing" sch_x=-210 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5787 N$22377 N$22379 N$22544 N$22546 "Waveguide Crossing" sch_x=-210 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5788 N$22381 N$22383 N$22548 N$22550 "Waveguide Crossing" sch_x=-210 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5789 N$22385 N$22387 N$22552 N$22554 "Waveguide Crossing" sch_x=-210 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5790 N$22389 N$22391 N$22556 N$22558 "Waveguide Crossing" sch_x=-210 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5791 N$22393 N$22395 N$22560 N$22562 "Waveguide Crossing" sch_x=-210 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5792 N$22397 N$22399 N$22564 N$22566 "Waveguide Crossing" sch_x=-210 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5793 N$22401 N$22403 N$22568 N$22570 "Waveguide Crossing" sch_x=-210 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5794 N$22405 N$22407 N$22572 N$22574 "Waveguide Crossing" sch_x=-210 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5795 N$22409 N$22411 N$22576 N$22578 "Waveguide Crossing" sch_x=-210 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5796 N$22413 N$22415 N$22580 N$22582 "Waveguide Crossing" sch_x=-210 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5797 N$22417 N$22419 N$22584 N$22586 "Waveguide Crossing" sch_x=-210 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5798 N$22421 N$22423 N$22588 N$22590 "Waveguide Crossing" sch_x=-210 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5799 N$22425 N$22427 N$22592 N$22594 "Waveguide Crossing" sch_x=-210 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5800 N$22429 N$22431 N$22596 N$22598 "Waveguide Crossing" sch_x=-210 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5801 N$22433 N$22435 N$22600 N$22602 "Waveguide Crossing" sch_x=-210 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5802 N$22437 N$22439 N$22604 N$22606 "Waveguide Crossing" sch_x=-210 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5803 N$22441 N$22443 N$22608 N$22610 "Waveguide Crossing" sch_x=-210 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5804 N$22445 N$22447 N$22612 N$22614 "Waveguide Crossing" sch_x=-210 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5805 N$22449 N$22451 N$22616 N$22618 "Waveguide Crossing" sch_x=-210 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5806 N$22453 N$22455 N$22620 N$22622 "Waveguide Crossing" sch_x=-210 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5807 N$22457 N$22459 N$22624 N$22626 "Waveguide Crossing" sch_x=-210 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5808 N$22461 N$22463 N$22628 N$22630 "Waveguide Crossing" sch_x=-210 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5809 N$22465 N$22467 N$22632 N$22634 "Waveguide Crossing" sch_x=-210 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5810 N$22469 N$22471 N$22636 N$22638 "Waveguide Crossing" sch_x=-210 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5811 N$22473 N$22475 N$22640 N$22642 "Waveguide Crossing" sch_x=-210 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5812 N$22477 N$22479 N$22644 N$22646 "Waveguide Crossing" sch_x=-210 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5813 N$22481 N$22483 N$22648 N$22650 "Waveguide Crossing" sch_x=-210 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5814 N$22485 N$22487 N$22652 N$22654 "Waveguide Crossing" sch_x=-210 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5815 N$22489 N$22491 N$22656 N$22658 "Waveguide Crossing" sch_x=-210 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5816 N$22493 N$22495 N$22660 N$22662 "Waveguide Crossing" sch_x=-210 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5817 N$22497 N$22499 N$22664 N$22666 "Waveguide Crossing" sch_x=-210 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5818 N$22501 N$22503 N$22668 N$22670 "Waveguide Crossing" sch_x=-210 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5819 N$22505 N$22507 N$22672 N$22674 "Waveguide Crossing" sch_x=-210 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5820 N$22509 N$22511 N$22676 N$22678 "Waveguide Crossing" sch_x=-210 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5821 N$22513 N$22515 N$22680 N$22682 "Waveguide Crossing" sch_x=-210 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5822 N$22517 N$22519 N$22684 N$22686 "Waveguide Crossing" sch_x=-210 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5823 N$22521 N$22523 N$22688 N$22690 "Waveguide Crossing" sch_x=-210 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5824 N$22525 N$22527 N$22692 N$22694 "Waveguide Crossing" sch_x=-210 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5825 N$22529 N$22531 N$22696 N$22698 "Waveguide Crossing" sch_x=-210 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5826 N$22533 N$22535 N$22700 N$22702 "Waveguide Crossing" sch_x=-210 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5827 N$22537 N$22539 N$22704 N$26193 "Waveguide Crossing" sch_x=-210 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5828 N$22541 N$22543 N$26029 N$22706 "Waveguide Crossing" sch_x=-208 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5829 N$22545 N$22547 N$22708 N$22710 "Waveguide Crossing" sch_x=-208 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5830 N$22549 N$22551 N$22712 N$22714 "Waveguide Crossing" sch_x=-208 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5831 N$22553 N$22555 N$22716 N$22718 "Waveguide Crossing" sch_x=-208 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5832 N$22557 N$22559 N$22720 N$22722 "Waveguide Crossing" sch_x=-208 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5833 N$22561 N$22563 N$22724 N$22726 "Waveguide Crossing" sch_x=-208 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5834 N$22565 N$22567 N$22728 N$22730 "Waveguide Crossing" sch_x=-208 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5835 N$22569 N$22571 N$22732 N$22734 "Waveguide Crossing" sch_x=-208 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5836 N$22573 N$22575 N$22736 N$22738 "Waveguide Crossing" sch_x=-208 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5837 N$22577 N$22579 N$22740 N$22742 "Waveguide Crossing" sch_x=-208 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5838 N$22581 N$22583 N$22744 N$22746 "Waveguide Crossing" sch_x=-208 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5839 N$22585 N$22587 N$22748 N$22750 "Waveguide Crossing" sch_x=-208 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5840 N$22589 N$22591 N$22752 N$22754 "Waveguide Crossing" sch_x=-208 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5841 N$22593 N$22595 N$22756 N$22758 "Waveguide Crossing" sch_x=-208 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5842 N$22597 N$22599 N$22760 N$22762 "Waveguide Crossing" sch_x=-208 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5843 N$22601 N$22603 N$22764 N$22766 "Waveguide Crossing" sch_x=-208 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5844 N$22605 N$22607 N$22768 N$22770 "Waveguide Crossing" sch_x=-208 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5845 N$22609 N$22611 N$22772 N$22774 "Waveguide Crossing" sch_x=-208 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5846 N$22613 N$22615 N$22776 N$22778 "Waveguide Crossing" sch_x=-208 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5847 N$22617 N$22619 N$22780 N$22782 "Waveguide Crossing" sch_x=-208 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5848 N$22621 N$22623 N$22784 N$22786 "Waveguide Crossing" sch_x=-208 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5849 N$22625 N$22627 N$22788 N$22790 "Waveguide Crossing" sch_x=-208 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5850 N$22629 N$22631 N$22792 N$22794 "Waveguide Crossing" sch_x=-208 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5851 N$22633 N$22635 N$22796 N$22798 "Waveguide Crossing" sch_x=-208 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5852 N$22637 N$22639 N$22800 N$22802 "Waveguide Crossing" sch_x=-208 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5853 N$22641 N$22643 N$22804 N$22806 "Waveguide Crossing" sch_x=-208 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5854 N$22645 N$22647 N$22808 N$22810 "Waveguide Crossing" sch_x=-208 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5855 N$22649 N$22651 N$22812 N$22814 "Waveguide Crossing" sch_x=-208 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5856 N$22653 N$22655 N$22816 N$22818 "Waveguide Crossing" sch_x=-208 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5857 N$22657 N$22659 N$22820 N$22822 "Waveguide Crossing" sch_x=-208 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5858 N$22661 N$22663 N$22824 N$22826 "Waveguide Crossing" sch_x=-208 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5859 N$22665 N$22667 N$22828 N$22830 "Waveguide Crossing" sch_x=-208 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5860 N$22669 N$22671 N$22832 N$22834 "Waveguide Crossing" sch_x=-208 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5861 N$22673 N$22675 N$22836 N$22838 "Waveguide Crossing" sch_x=-208 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5862 N$22677 N$22679 N$22840 N$22842 "Waveguide Crossing" sch_x=-208 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5863 N$22681 N$22683 N$22844 N$22846 "Waveguide Crossing" sch_x=-208 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5864 N$22685 N$22687 N$22848 N$22850 "Waveguide Crossing" sch_x=-208 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5865 N$22689 N$22691 N$22852 N$22854 "Waveguide Crossing" sch_x=-208 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5866 N$22693 N$22695 N$22856 N$22858 "Waveguide Crossing" sch_x=-208 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5867 N$22697 N$22699 N$22860 N$22862 "Waveguide Crossing" sch_x=-208 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5868 N$22701 N$22703 N$22864 N$26191 "Waveguide Crossing" sch_x=-208 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5869 N$22705 N$22707 N$26031 N$22866 "Waveguide Crossing" sch_x=-206 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5870 N$22709 N$22711 N$22868 N$22870 "Waveguide Crossing" sch_x=-206 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5871 N$22713 N$22715 N$22872 N$22874 "Waveguide Crossing" sch_x=-206 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5872 N$22717 N$22719 N$22876 N$22878 "Waveguide Crossing" sch_x=-206 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5873 N$22721 N$22723 N$22880 N$22882 "Waveguide Crossing" sch_x=-206 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5874 N$22725 N$22727 N$22884 N$22886 "Waveguide Crossing" sch_x=-206 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5875 N$22729 N$22731 N$22888 N$22890 "Waveguide Crossing" sch_x=-206 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5876 N$22733 N$22735 N$22892 N$22894 "Waveguide Crossing" sch_x=-206 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5877 N$22737 N$22739 N$22896 N$22898 "Waveguide Crossing" sch_x=-206 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5878 N$22741 N$22743 N$22900 N$22902 "Waveguide Crossing" sch_x=-206 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5879 N$22745 N$22747 N$22904 N$22906 "Waveguide Crossing" sch_x=-206 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5880 N$22749 N$22751 N$22908 N$22910 "Waveguide Crossing" sch_x=-206 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5881 N$22753 N$22755 N$22912 N$22914 "Waveguide Crossing" sch_x=-206 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5882 N$22757 N$22759 N$22916 N$22918 "Waveguide Crossing" sch_x=-206 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5883 N$22761 N$22763 N$22920 N$22922 "Waveguide Crossing" sch_x=-206 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5884 N$22765 N$22767 N$22924 N$22926 "Waveguide Crossing" sch_x=-206 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5885 N$22769 N$22771 N$22928 N$22930 "Waveguide Crossing" sch_x=-206 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5886 N$22773 N$22775 N$22932 N$22934 "Waveguide Crossing" sch_x=-206 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5887 N$22777 N$22779 N$22936 N$22938 "Waveguide Crossing" sch_x=-206 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5888 N$22781 N$22783 N$22940 N$22942 "Waveguide Crossing" sch_x=-206 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5889 N$22785 N$22787 N$22944 N$22946 "Waveguide Crossing" sch_x=-206 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5890 N$22789 N$22791 N$22948 N$22950 "Waveguide Crossing" sch_x=-206 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5891 N$22793 N$22795 N$22952 N$22954 "Waveguide Crossing" sch_x=-206 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5892 N$22797 N$22799 N$22956 N$22958 "Waveguide Crossing" sch_x=-206 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5893 N$22801 N$22803 N$22960 N$22962 "Waveguide Crossing" sch_x=-206 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5894 N$22805 N$22807 N$22964 N$22966 "Waveguide Crossing" sch_x=-206 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5895 N$22809 N$22811 N$22968 N$22970 "Waveguide Crossing" sch_x=-206 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5896 N$22813 N$22815 N$22972 N$22974 "Waveguide Crossing" sch_x=-206 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5897 N$22817 N$22819 N$22976 N$22978 "Waveguide Crossing" sch_x=-206 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5898 N$22821 N$22823 N$22980 N$22982 "Waveguide Crossing" sch_x=-206 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5899 N$22825 N$22827 N$22984 N$22986 "Waveguide Crossing" sch_x=-206 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5900 N$22829 N$22831 N$22988 N$22990 "Waveguide Crossing" sch_x=-206 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5901 N$22833 N$22835 N$22992 N$22994 "Waveguide Crossing" sch_x=-206 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5902 N$22837 N$22839 N$22996 N$22998 "Waveguide Crossing" sch_x=-206 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5903 N$22841 N$22843 N$23000 N$23002 "Waveguide Crossing" sch_x=-206 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5904 N$22845 N$22847 N$23004 N$23006 "Waveguide Crossing" sch_x=-206 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5905 N$22849 N$22851 N$23008 N$23010 "Waveguide Crossing" sch_x=-206 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5906 N$22853 N$22855 N$23012 N$23014 "Waveguide Crossing" sch_x=-206 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5907 N$22857 N$22859 N$23016 N$23018 "Waveguide Crossing" sch_x=-206 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5908 N$22861 N$22863 N$23020 N$26189 "Waveguide Crossing" sch_x=-206 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5909 N$22865 N$22867 N$26033 N$23022 "Waveguide Crossing" sch_x=-204 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5910 N$22869 N$22871 N$23024 N$23026 "Waveguide Crossing" sch_x=-204 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5911 N$22873 N$22875 N$23028 N$23030 "Waveguide Crossing" sch_x=-204 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5912 N$22877 N$22879 N$23032 N$23034 "Waveguide Crossing" sch_x=-204 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5913 N$22881 N$22883 N$23036 N$23038 "Waveguide Crossing" sch_x=-204 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5914 N$22885 N$22887 N$23040 N$23042 "Waveguide Crossing" sch_x=-204 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5915 N$22889 N$22891 N$23044 N$23046 "Waveguide Crossing" sch_x=-204 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5916 N$22893 N$22895 N$23048 N$23050 "Waveguide Crossing" sch_x=-204 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5917 N$22897 N$22899 N$23052 N$23054 "Waveguide Crossing" sch_x=-204 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5918 N$22901 N$22903 N$23056 N$23058 "Waveguide Crossing" sch_x=-204 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5919 N$22905 N$22907 N$23060 N$23062 "Waveguide Crossing" sch_x=-204 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5920 N$22909 N$22911 N$23064 N$23066 "Waveguide Crossing" sch_x=-204 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5921 N$22913 N$22915 N$23068 N$23070 "Waveguide Crossing" sch_x=-204 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5922 N$22917 N$22919 N$23072 N$23074 "Waveguide Crossing" sch_x=-204 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5923 N$22921 N$22923 N$23076 N$23078 "Waveguide Crossing" sch_x=-204 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5924 N$22925 N$22927 N$23080 N$23082 "Waveguide Crossing" sch_x=-204 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5925 N$22929 N$22931 N$23084 N$23086 "Waveguide Crossing" sch_x=-204 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5926 N$22933 N$22935 N$23088 N$23090 "Waveguide Crossing" sch_x=-204 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5927 N$22937 N$22939 N$23092 N$23094 "Waveguide Crossing" sch_x=-204 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5928 N$22941 N$22943 N$23096 N$23098 "Waveguide Crossing" sch_x=-204 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5929 N$22945 N$22947 N$23100 N$23102 "Waveguide Crossing" sch_x=-204 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5930 N$22949 N$22951 N$23104 N$23106 "Waveguide Crossing" sch_x=-204 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5931 N$22953 N$22955 N$23108 N$23110 "Waveguide Crossing" sch_x=-204 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5932 N$22957 N$22959 N$23112 N$23114 "Waveguide Crossing" sch_x=-204 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5933 N$22961 N$22963 N$23116 N$23118 "Waveguide Crossing" sch_x=-204 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5934 N$22965 N$22967 N$23120 N$23122 "Waveguide Crossing" sch_x=-204 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5935 N$22969 N$22971 N$23124 N$23126 "Waveguide Crossing" sch_x=-204 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5936 N$22973 N$22975 N$23128 N$23130 "Waveguide Crossing" sch_x=-204 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5937 N$22977 N$22979 N$23132 N$23134 "Waveguide Crossing" sch_x=-204 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5938 N$22981 N$22983 N$23136 N$23138 "Waveguide Crossing" sch_x=-204 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5939 N$22985 N$22987 N$23140 N$23142 "Waveguide Crossing" sch_x=-204 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5940 N$22989 N$22991 N$23144 N$23146 "Waveguide Crossing" sch_x=-204 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5941 N$22993 N$22995 N$23148 N$23150 "Waveguide Crossing" sch_x=-204 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5942 N$22997 N$22999 N$23152 N$23154 "Waveguide Crossing" sch_x=-204 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5943 N$23001 N$23003 N$23156 N$23158 "Waveguide Crossing" sch_x=-204 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5944 N$23005 N$23007 N$23160 N$23162 "Waveguide Crossing" sch_x=-204 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5945 N$23009 N$23011 N$23164 N$23166 "Waveguide Crossing" sch_x=-204 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5946 N$23013 N$23015 N$23168 N$23170 "Waveguide Crossing" sch_x=-204 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5947 N$23017 N$23019 N$23172 N$26187 "Waveguide Crossing" sch_x=-204 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5948 N$23021 N$23023 N$26035 N$23174 "Waveguide Crossing" sch_x=-202 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5949 N$23025 N$23027 N$23176 N$23178 "Waveguide Crossing" sch_x=-202 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5950 N$23029 N$23031 N$23180 N$23182 "Waveguide Crossing" sch_x=-202 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5951 N$23033 N$23035 N$23184 N$23186 "Waveguide Crossing" sch_x=-202 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5952 N$23037 N$23039 N$23188 N$23190 "Waveguide Crossing" sch_x=-202 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5953 N$23041 N$23043 N$23192 N$23194 "Waveguide Crossing" sch_x=-202 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5954 N$23045 N$23047 N$23196 N$23198 "Waveguide Crossing" sch_x=-202 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5955 N$23049 N$23051 N$23200 N$23202 "Waveguide Crossing" sch_x=-202 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5956 N$23053 N$23055 N$23204 N$23206 "Waveguide Crossing" sch_x=-202 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5957 N$23057 N$23059 N$23208 N$23210 "Waveguide Crossing" sch_x=-202 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5958 N$23061 N$23063 N$23212 N$23214 "Waveguide Crossing" sch_x=-202 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5959 N$23065 N$23067 N$23216 N$23218 "Waveguide Crossing" sch_x=-202 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5960 N$23069 N$23071 N$23220 N$23222 "Waveguide Crossing" sch_x=-202 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5961 N$23073 N$23075 N$23224 N$23226 "Waveguide Crossing" sch_x=-202 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5962 N$23077 N$23079 N$23228 N$23230 "Waveguide Crossing" sch_x=-202 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5963 N$23081 N$23083 N$23232 N$23234 "Waveguide Crossing" sch_x=-202 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5964 N$23085 N$23087 N$23236 N$23238 "Waveguide Crossing" sch_x=-202 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5965 N$23089 N$23091 N$23240 N$23242 "Waveguide Crossing" sch_x=-202 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5966 N$23093 N$23095 N$23244 N$23246 "Waveguide Crossing" sch_x=-202 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5967 N$23097 N$23099 N$23248 N$23250 "Waveguide Crossing" sch_x=-202 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5968 N$23101 N$23103 N$23252 N$23254 "Waveguide Crossing" sch_x=-202 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5969 N$23105 N$23107 N$23256 N$23258 "Waveguide Crossing" sch_x=-202 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5970 N$23109 N$23111 N$23260 N$23262 "Waveguide Crossing" sch_x=-202 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5971 N$23113 N$23115 N$23264 N$23266 "Waveguide Crossing" sch_x=-202 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5972 N$23117 N$23119 N$23268 N$23270 "Waveguide Crossing" sch_x=-202 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5973 N$23121 N$23123 N$23272 N$23274 "Waveguide Crossing" sch_x=-202 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5974 N$23125 N$23127 N$23276 N$23278 "Waveguide Crossing" sch_x=-202 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5975 N$23129 N$23131 N$23280 N$23282 "Waveguide Crossing" sch_x=-202 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5976 N$23133 N$23135 N$23284 N$23286 "Waveguide Crossing" sch_x=-202 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5977 N$23137 N$23139 N$23288 N$23290 "Waveguide Crossing" sch_x=-202 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5978 N$23141 N$23143 N$23292 N$23294 "Waveguide Crossing" sch_x=-202 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5979 N$23145 N$23147 N$23296 N$23298 "Waveguide Crossing" sch_x=-202 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5980 N$23149 N$23151 N$23300 N$23302 "Waveguide Crossing" sch_x=-202 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5981 N$23153 N$23155 N$23304 N$23306 "Waveguide Crossing" sch_x=-202 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5982 N$23157 N$23159 N$23308 N$23310 "Waveguide Crossing" sch_x=-202 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5983 N$23161 N$23163 N$23312 N$23314 "Waveguide Crossing" sch_x=-202 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5984 N$23165 N$23167 N$23316 N$23318 "Waveguide Crossing" sch_x=-202 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5985 N$23169 N$23171 N$23320 N$26185 "Waveguide Crossing" sch_x=-202 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5986 N$23173 N$23175 N$26037 N$23322 "Waveguide Crossing" sch_x=-200 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5987 N$23177 N$23179 N$23324 N$23326 "Waveguide Crossing" sch_x=-200 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5988 N$23181 N$23183 N$23328 N$23330 "Waveguide Crossing" sch_x=-200 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5989 N$23185 N$23187 N$23332 N$23334 "Waveguide Crossing" sch_x=-200 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5990 N$23189 N$23191 N$23336 N$23338 "Waveguide Crossing" sch_x=-200 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5991 N$23193 N$23195 N$23340 N$23342 "Waveguide Crossing" sch_x=-200 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5992 N$23197 N$23199 N$23344 N$23346 "Waveguide Crossing" sch_x=-200 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5993 N$23201 N$23203 N$23348 N$23350 "Waveguide Crossing" sch_x=-200 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5994 N$23205 N$23207 N$23352 N$23354 "Waveguide Crossing" sch_x=-200 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5995 N$23209 N$23211 N$23356 N$23358 "Waveguide Crossing" sch_x=-200 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5996 N$23213 N$23215 N$23360 N$23362 "Waveguide Crossing" sch_x=-200 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5997 N$23217 N$23219 N$23364 N$23366 "Waveguide Crossing" sch_x=-200 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5998 N$23221 N$23223 N$23368 N$23370 "Waveguide Crossing" sch_x=-200 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C5999 N$23225 N$23227 N$23372 N$23374 "Waveguide Crossing" sch_x=-200 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6000 N$23229 N$23231 N$23376 N$23378 "Waveguide Crossing" sch_x=-200 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6001 N$23233 N$23235 N$23380 N$23382 "Waveguide Crossing" sch_x=-200 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6002 N$23237 N$23239 N$23384 N$23386 "Waveguide Crossing" sch_x=-200 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6003 N$23241 N$23243 N$23388 N$23390 "Waveguide Crossing" sch_x=-200 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6004 N$23245 N$23247 N$23392 N$23394 "Waveguide Crossing" sch_x=-200 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6005 N$23249 N$23251 N$23396 N$23398 "Waveguide Crossing" sch_x=-200 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6006 N$23253 N$23255 N$23400 N$23402 "Waveguide Crossing" sch_x=-200 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6007 N$23257 N$23259 N$23404 N$23406 "Waveguide Crossing" sch_x=-200 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6008 N$23261 N$23263 N$23408 N$23410 "Waveguide Crossing" sch_x=-200 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6009 N$23265 N$23267 N$23412 N$23414 "Waveguide Crossing" sch_x=-200 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6010 N$23269 N$23271 N$23416 N$23418 "Waveguide Crossing" sch_x=-200 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6011 N$23273 N$23275 N$23420 N$23422 "Waveguide Crossing" sch_x=-200 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6012 N$23277 N$23279 N$23424 N$23426 "Waveguide Crossing" sch_x=-200 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6013 N$23281 N$23283 N$23428 N$23430 "Waveguide Crossing" sch_x=-200 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6014 N$23285 N$23287 N$23432 N$23434 "Waveguide Crossing" sch_x=-200 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6015 N$23289 N$23291 N$23436 N$23438 "Waveguide Crossing" sch_x=-200 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6016 N$23293 N$23295 N$23440 N$23442 "Waveguide Crossing" sch_x=-200 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6017 N$23297 N$23299 N$23444 N$23446 "Waveguide Crossing" sch_x=-200 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6018 N$23301 N$23303 N$23448 N$23450 "Waveguide Crossing" sch_x=-200 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6019 N$23305 N$23307 N$23452 N$23454 "Waveguide Crossing" sch_x=-200 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6020 N$23309 N$23311 N$23456 N$23458 "Waveguide Crossing" sch_x=-200 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6021 N$23313 N$23315 N$23460 N$23462 "Waveguide Crossing" sch_x=-200 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6022 N$23317 N$23319 N$23464 N$26183 "Waveguide Crossing" sch_x=-200 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6023 N$23321 N$23323 N$26039 N$23466 "Waveguide Crossing" sch_x=-198 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6024 N$23325 N$23327 N$23468 N$23470 "Waveguide Crossing" sch_x=-198 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6025 N$23329 N$23331 N$23472 N$23474 "Waveguide Crossing" sch_x=-198 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6026 N$23333 N$23335 N$23476 N$23478 "Waveguide Crossing" sch_x=-198 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6027 N$23337 N$23339 N$23480 N$23482 "Waveguide Crossing" sch_x=-198 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6028 N$23341 N$23343 N$23484 N$23486 "Waveguide Crossing" sch_x=-198 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6029 N$23345 N$23347 N$23488 N$23490 "Waveguide Crossing" sch_x=-198 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6030 N$23349 N$23351 N$23492 N$23494 "Waveguide Crossing" sch_x=-198 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6031 N$23353 N$23355 N$23496 N$23498 "Waveguide Crossing" sch_x=-198 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6032 N$23357 N$23359 N$23500 N$23502 "Waveguide Crossing" sch_x=-198 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6033 N$23361 N$23363 N$23504 N$23506 "Waveguide Crossing" sch_x=-198 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6034 N$23365 N$23367 N$23508 N$23510 "Waveguide Crossing" sch_x=-198 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6035 N$23369 N$23371 N$23512 N$23514 "Waveguide Crossing" sch_x=-198 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6036 N$23373 N$23375 N$23516 N$23518 "Waveguide Crossing" sch_x=-198 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6037 N$23377 N$23379 N$23520 N$23522 "Waveguide Crossing" sch_x=-198 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6038 N$23381 N$23383 N$23524 N$23526 "Waveguide Crossing" sch_x=-198 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6039 N$23385 N$23387 N$23528 N$23530 "Waveguide Crossing" sch_x=-198 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6040 N$23389 N$23391 N$23532 N$23534 "Waveguide Crossing" sch_x=-198 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6041 N$23393 N$23395 N$23536 N$23538 "Waveguide Crossing" sch_x=-198 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6042 N$23397 N$23399 N$23540 N$23542 "Waveguide Crossing" sch_x=-198 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6043 N$23401 N$23403 N$23544 N$23546 "Waveguide Crossing" sch_x=-198 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6044 N$23405 N$23407 N$23548 N$23550 "Waveguide Crossing" sch_x=-198 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6045 N$23409 N$23411 N$23552 N$23554 "Waveguide Crossing" sch_x=-198 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6046 N$23413 N$23415 N$23556 N$23558 "Waveguide Crossing" sch_x=-198 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6047 N$23417 N$23419 N$23560 N$23562 "Waveguide Crossing" sch_x=-198 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6048 N$23421 N$23423 N$23564 N$23566 "Waveguide Crossing" sch_x=-198 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6049 N$23425 N$23427 N$23568 N$23570 "Waveguide Crossing" sch_x=-198 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6050 N$23429 N$23431 N$23572 N$23574 "Waveguide Crossing" sch_x=-198 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6051 N$23433 N$23435 N$23576 N$23578 "Waveguide Crossing" sch_x=-198 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6052 N$23437 N$23439 N$23580 N$23582 "Waveguide Crossing" sch_x=-198 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6053 N$23441 N$23443 N$23584 N$23586 "Waveguide Crossing" sch_x=-198 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6054 N$23445 N$23447 N$23588 N$23590 "Waveguide Crossing" sch_x=-198 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6055 N$23449 N$23451 N$23592 N$23594 "Waveguide Crossing" sch_x=-198 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6056 N$23453 N$23455 N$23596 N$23598 "Waveguide Crossing" sch_x=-198 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6057 N$23457 N$23459 N$23600 N$23602 "Waveguide Crossing" sch_x=-198 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6058 N$23461 N$23463 N$23604 N$26181 "Waveguide Crossing" sch_x=-198 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6059 N$23465 N$23467 N$26041 N$23606 "Waveguide Crossing" sch_x=-196 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6060 N$23469 N$23471 N$23608 N$23610 "Waveguide Crossing" sch_x=-196 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6061 N$23473 N$23475 N$23612 N$23614 "Waveguide Crossing" sch_x=-196 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6062 N$23477 N$23479 N$23616 N$23618 "Waveguide Crossing" sch_x=-196 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6063 N$23481 N$23483 N$23620 N$23622 "Waveguide Crossing" sch_x=-196 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6064 N$23485 N$23487 N$23624 N$23626 "Waveguide Crossing" sch_x=-196 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6065 N$23489 N$23491 N$23628 N$23630 "Waveguide Crossing" sch_x=-196 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6066 N$23493 N$23495 N$23632 N$23634 "Waveguide Crossing" sch_x=-196 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6067 N$23497 N$23499 N$23636 N$23638 "Waveguide Crossing" sch_x=-196 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6068 N$23501 N$23503 N$23640 N$23642 "Waveguide Crossing" sch_x=-196 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6069 N$23505 N$23507 N$23644 N$23646 "Waveguide Crossing" sch_x=-196 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6070 N$23509 N$23511 N$23648 N$23650 "Waveguide Crossing" sch_x=-196 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6071 N$23513 N$23515 N$23652 N$23654 "Waveguide Crossing" sch_x=-196 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6072 N$23517 N$23519 N$23656 N$23658 "Waveguide Crossing" sch_x=-196 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6073 N$23521 N$23523 N$23660 N$23662 "Waveguide Crossing" sch_x=-196 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6074 N$23525 N$23527 N$23664 N$23666 "Waveguide Crossing" sch_x=-196 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6075 N$23529 N$23531 N$23668 N$23670 "Waveguide Crossing" sch_x=-196 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6076 N$23533 N$23535 N$23672 N$23674 "Waveguide Crossing" sch_x=-196 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6077 N$23537 N$23539 N$23676 N$23678 "Waveguide Crossing" sch_x=-196 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6078 N$23541 N$23543 N$23680 N$23682 "Waveguide Crossing" sch_x=-196 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6079 N$23545 N$23547 N$23684 N$23686 "Waveguide Crossing" sch_x=-196 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6080 N$23549 N$23551 N$23688 N$23690 "Waveguide Crossing" sch_x=-196 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6081 N$23553 N$23555 N$23692 N$23694 "Waveguide Crossing" sch_x=-196 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6082 N$23557 N$23559 N$23696 N$23698 "Waveguide Crossing" sch_x=-196 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6083 N$23561 N$23563 N$23700 N$23702 "Waveguide Crossing" sch_x=-196 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6084 N$23565 N$23567 N$23704 N$23706 "Waveguide Crossing" sch_x=-196 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6085 N$23569 N$23571 N$23708 N$23710 "Waveguide Crossing" sch_x=-196 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6086 N$23573 N$23575 N$23712 N$23714 "Waveguide Crossing" sch_x=-196 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6087 N$23577 N$23579 N$23716 N$23718 "Waveguide Crossing" sch_x=-196 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6088 N$23581 N$23583 N$23720 N$23722 "Waveguide Crossing" sch_x=-196 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6089 N$23585 N$23587 N$23724 N$23726 "Waveguide Crossing" sch_x=-196 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6090 N$23589 N$23591 N$23728 N$23730 "Waveguide Crossing" sch_x=-196 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6091 N$23593 N$23595 N$23732 N$23734 "Waveguide Crossing" sch_x=-196 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6092 N$23597 N$23599 N$23736 N$23738 "Waveguide Crossing" sch_x=-196 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6093 N$23601 N$23603 N$23740 N$26179 "Waveguide Crossing" sch_x=-196 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6094 N$23605 N$23607 N$26043 N$23742 "Waveguide Crossing" sch_x=-194 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6095 N$23609 N$23611 N$23744 N$23746 "Waveguide Crossing" sch_x=-194 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6096 N$23613 N$23615 N$23748 N$23750 "Waveguide Crossing" sch_x=-194 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6097 N$23617 N$23619 N$23752 N$23754 "Waveguide Crossing" sch_x=-194 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6098 N$23621 N$23623 N$23756 N$23758 "Waveguide Crossing" sch_x=-194 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6099 N$23625 N$23627 N$23760 N$23762 "Waveguide Crossing" sch_x=-194 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6100 N$23629 N$23631 N$23764 N$23766 "Waveguide Crossing" sch_x=-194 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6101 N$23633 N$23635 N$23768 N$23770 "Waveguide Crossing" sch_x=-194 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6102 N$23637 N$23639 N$23772 N$23774 "Waveguide Crossing" sch_x=-194 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6103 N$23641 N$23643 N$23776 N$23778 "Waveguide Crossing" sch_x=-194 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6104 N$23645 N$23647 N$23780 N$23782 "Waveguide Crossing" sch_x=-194 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6105 N$23649 N$23651 N$23784 N$23786 "Waveguide Crossing" sch_x=-194 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6106 N$23653 N$23655 N$23788 N$23790 "Waveguide Crossing" sch_x=-194 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6107 N$23657 N$23659 N$23792 N$23794 "Waveguide Crossing" sch_x=-194 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6108 N$23661 N$23663 N$23796 N$23798 "Waveguide Crossing" sch_x=-194 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6109 N$23665 N$23667 N$23800 N$23802 "Waveguide Crossing" sch_x=-194 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6110 N$23669 N$23671 N$23804 N$23806 "Waveguide Crossing" sch_x=-194 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6111 N$23673 N$23675 N$23808 N$23810 "Waveguide Crossing" sch_x=-194 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6112 N$23677 N$23679 N$23812 N$23814 "Waveguide Crossing" sch_x=-194 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6113 N$23681 N$23683 N$23816 N$23818 "Waveguide Crossing" sch_x=-194 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6114 N$23685 N$23687 N$23820 N$23822 "Waveguide Crossing" sch_x=-194 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6115 N$23689 N$23691 N$23824 N$23826 "Waveguide Crossing" sch_x=-194 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6116 N$23693 N$23695 N$23828 N$23830 "Waveguide Crossing" sch_x=-194 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6117 N$23697 N$23699 N$23832 N$23834 "Waveguide Crossing" sch_x=-194 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6118 N$23701 N$23703 N$23836 N$23838 "Waveguide Crossing" sch_x=-194 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6119 N$23705 N$23707 N$23840 N$23842 "Waveguide Crossing" sch_x=-194 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6120 N$23709 N$23711 N$23844 N$23846 "Waveguide Crossing" sch_x=-194 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6121 N$23713 N$23715 N$23848 N$23850 "Waveguide Crossing" sch_x=-194 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6122 N$23717 N$23719 N$23852 N$23854 "Waveguide Crossing" sch_x=-194 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6123 N$23721 N$23723 N$23856 N$23858 "Waveguide Crossing" sch_x=-194 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6124 N$23725 N$23727 N$23860 N$23862 "Waveguide Crossing" sch_x=-194 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6125 N$23729 N$23731 N$23864 N$23866 "Waveguide Crossing" sch_x=-194 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6126 N$23733 N$23735 N$23868 N$23870 "Waveguide Crossing" sch_x=-194 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6127 N$23737 N$23739 N$23872 N$26177 "Waveguide Crossing" sch_x=-194 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6128 N$23741 N$23743 N$26045 N$23874 "Waveguide Crossing" sch_x=-192 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6129 N$23745 N$23747 N$23876 N$23878 "Waveguide Crossing" sch_x=-192 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6130 N$23749 N$23751 N$23880 N$23882 "Waveguide Crossing" sch_x=-192 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6131 N$23753 N$23755 N$23884 N$23886 "Waveguide Crossing" sch_x=-192 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6132 N$23757 N$23759 N$23888 N$23890 "Waveguide Crossing" sch_x=-192 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6133 N$23761 N$23763 N$23892 N$23894 "Waveguide Crossing" sch_x=-192 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6134 N$23765 N$23767 N$23896 N$23898 "Waveguide Crossing" sch_x=-192 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6135 N$23769 N$23771 N$23900 N$23902 "Waveguide Crossing" sch_x=-192 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6136 N$23773 N$23775 N$23904 N$23906 "Waveguide Crossing" sch_x=-192 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6137 N$23777 N$23779 N$23908 N$23910 "Waveguide Crossing" sch_x=-192 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6138 N$23781 N$23783 N$23912 N$23914 "Waveguide Crossing" sch_x=-192 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6139 N$23785 N$23787 N$23916 N$23918 "Waveguide Crossing" sch_x=-192 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6140 N$23789 N$23791 N$23920 N$23922 "Waveguide Crossing" sch_x=-192 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6141 N$23793 N$23795 N$23924 N$23926 "Waveguide Crossing" sch_x=-192 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6142 N$23797 N$23799 N$23928 N$23930 "Waveguide Crossing" sch_x=-192 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6143 N$23801 N$23803 N$23932 N$23934 "Waveguide Crossing" sch_x=-192 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6144 N$23805 N$23807 N$23936 N$23938 "Waveguide Crossing" sch_x=-192 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6145 N$23809 N$23811 N$23940 N$23942 "Waveguide Crossing" sch_x=-192 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6146 N$23813 N$23815 N$23944 N$23946 "Waveguide Crossing" sch_x=-192 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6147 N$23817 N$23819 N$23948 N$23950 "Waveguide Crossing" sch_x=-192 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6148 N$23821 N$23823 N$23952 N$23954 "Waveguide Crossing" sch_x=-192 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6149 N$23825 N$23827 N$23956 N$23958 "Waveguide Crossing" sch_x=-192 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6150 N$23829 N$23831 N$23960 N$23962 "Waveguide Crossing" sch_x=-192 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6151 N$23833 N$23835 N$23964 N$23966 "Waveguide Crossing" sch_x=-192 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6152 N$23837 N$23839 N$23968 N$23970 "Waveguide Crossing" sch_x=-192 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6153 N$23841 N$23843 N$23972 N$23974 "Waveguide Crossing" sch_x=-192 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6154 N$23845 N$23847 N$23976 N$23978 "Waveguide Crossing" sch_x=-192 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6155 N$23849 N$23851 N$23980 N$23982 "Waveguide Crossing" sch_x=-192 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6156 N$23853 N$23855 N$23984 N$23986 "Waveguide Crossing" sch_x=-192 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6157 N$23857 N$23859 N$23988 N$23990 "Waveguide Crossing" sch_x=-192 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6158 N$23861 N$23863 N$23992 N$23994 "Waveguide Crossing" sch_x=-192 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6159 N$23865 N$23867 N$23996 N$23998 "Waveguide Crossing" sch_x=-192 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6160 N$23869 N$23871 N$24000 N$26175 "Waveguide Crossing" sch_x=-192 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6161 N$23873 N$23875 N$26047 N$24002 "Waveguide Crossing" sch_x=-190 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6162 N$23877 N$23879 N$24004 N$24006 "Waveguide Crossing" sch_x=-190 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6163 N$23881 N$23883 N$24008 N$24010 "Waveguide Crossing" sch_x=-190 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6164 N$23885 N$23887 N$24012 N$24014 "Waveguide Crossing" sch_x=-190 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6165 N$23889 N$23891 N$24016 N$24018 "Waveguide Crossing" sch_x=-190 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6166 N$23893 N$23895 N$24020 N$24022 "Waveguide Crossing" sch_x=-190 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6167 N$23897 N$23899 N$24024 N$24026 "Waveguide Crossing" sch_x=-190 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6168 N$23901 N$23903 N$24028 N$24030 "Waveguide Crossing" sch_x=-190 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6169 N$23905 N$23907 N$24032 N$24034 "Waveguide Crossing" sch_x=-190 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6170 N$23909 N$23911 N$24036 N$24038 "Waveguide Crossing" sch_x=-190 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6171 N$23913 N$23915 N$24040 N$24042 "Waveguide Crossing" sch_x=-190 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6172 N$23917 N$23919 N$24044 N$24046 "Waveguide Crossing" sch_x=-190 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6173 N$23921 N$23923 N$24048 N$24050 "Waveguide Crossing" sch_x=-190 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6174 N$23925 N$23927 N$24052 N$24054 "Waveguide Crossing" sch_x=-190 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6175 N$23929 N$23931 N$24056 N$24058 "Waveguide Crossing" sch_x=-190 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6176 N$23933 N$23935 N$24060 N$24062 "Waveguide Crossing" sch_x=-190 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6177 N$23937 N$23939 N$24064 N$24066 "Waveguide Crossing" sch_x=-190 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6178 N$23941 N$23943 N$24068 N$24070 "Waveguide Crossing" sch_x=-190 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6179 N$23945 N$23947 N$24072 N$24074 "Waveguide Crossing" sch_x=-190 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6180 N$23949 N$23951 N$24076 N$24078 "Waveguide Crossing" sch_x=-190 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6181 N$23953 N$23955 N$24080 N$24082 "Waveguide Crossing" sch_x=-190 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6182 N$23957 N$23959 N$24084 N$24086 "Waveguide Crossing" sch_x=-190 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6183 N$23961 N$23963 N$24088 N$24090 "Waveguide Crossing" sch_x=-190 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6184 N$23965 N$23967 N$24092 N$24094 "Waveguide Crossing" sch_x=-190 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6185 N$23969 N$23971 N$24096 N$24098 "Waveguide Crossing" sch_x=-190 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6186 N$23973 N$23975 N$24100 N$24102 "Waveguide Crossing" sch_x=-190 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6187 N$23977 N$23979 N$24104 N$24106 "Waveguide Crossing" sch_x=-190 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6188 N$23981 N$23983 N$24108 N$24110 "Waveguide Crossing" sch_x=-190 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6189 N$23985 N$23987 N$24112 N$24114 "Waveguide Crossing" sch_x=-190 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6190 N$23989 N$23991 N$24116 N$24118 "Waveguide Crossing" sch_x=-190 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6191 N$23993 N$23995 N$24120 N$24122 "Waveguide Crossing" sch_x=-190 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6192 N$23997 N$23999 N$24124 N$26173 "Waveguide Crossing" sch_x=-190 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6193 N$24001 N$24003 N$26049 N$24126 "Waveguide Crossing" sch_x=-188 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6194 N$24005 N$24007 N$24128 N$24130 "Waveguide Crossing" sch_x=-188 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6195 N$24009 N$24011 N$24132 N$24134 "Waveguide Crossing" sch_x=-188 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6196 N$24013 N$24015 N$24136 N$24138 "Waveguide Crossing" sch_x=-188 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6197 N$24017 N$24019 N$24140 N$24142 "Waveguide Crossing" sch_x=-188 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6198 N$24021 N$24023 N$24144 N$24146 "Waveguide Crossing" sch_x=-188 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6199 N$24025 N$24027 N$24148 N$24150 "Waveguide Crossing" sch_x=-188 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6200 N$24029 N$24031 N$24152 N$24154 "Waveguide Crossing" sch_x=-188 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6201 N$24033 N$24035 N$24156 N$24158 "Waveguide Crossing" sch_x=-188 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6202 N$24037 N$24039 N$24160 N$24162 "Waveguide Crossing" sch_x=-188 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6203 N$24041 N$24043 N$24164 N$24166 "Waveguide Crossing" sch_x=-188 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6204 N$24045 N$24047 N$24168 N$24170 "Waveguide Crossing" sch_x=-188 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6205 N$24049 N$24051 N$24172 N$24174 "Waveguide Crossing" sch_x=-188 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6206 N$24053 N$24055 N$24176 N$24178 "Waveguide Crossing" sch_x=-188 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6207 N$24057 N$24059 N$24180 N$24182 "Waveguide Crossing" sch_x=-188 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6208 N$24061 N$24063 N$24184 N$24186 "Waveguide Crossing" sch_x=-188 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6209 N$24065 N$24067 N$24188 N$24190 "Waveguide Crossing" sch_x=-188 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6210 N$24069 N$24071 N$24192 N$24194 "Waveguide Crossing" sch_x=-188 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6211 N$24073 N$24075 N$24196 N$24198 "Waveguide Crossing" sch_x=-188 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6212 N$24077 N$24079 N$24200 N$24202 "Waveguide Crossing" sch_x=-188 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6213 N$24081 N$24083 N$24204 N$24206 "Waveguide Crossing" sch_x=-188 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6214 N$24085 N$24087 N$24208 N$24210 "Waveguide Crossing" sch_x=-188 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6215 N$24089 N$24091 N$24212 N$24214 "Waveguide Crossing" sch_x=-188 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6216 N$24093 N$24095 N$24216 N$24218 "Waveguide Crossing" sch_x=-188 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6217 N$24097 N$24099 N$24220 N$24222 "Waveguide Crossing" sch_x=-188 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6218 N$24101 N$24103 N$24224 N$24226 "Waveguide Crossing" sch_x=-188 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6219 N$24105 N$24107 N$24228 N$24230 "Waveguide Crossing" sch_x=-188 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6220 N$24109 N$24111 N$24232 N$24234 "Waveguide Crossing" sch_x=-188 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6221 N$24113 N$24115 N$24236 N$24238 "Waveguide Crossing" sch_x=-188 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6222 N$24117 N$24119 N$24240 N$24242 "Waveguide Crossing" sch_x=-188 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6223 N$24121 N$24123 N$24244 N$26171 "Waveguide Crossing" sch_x=-188 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6224 N$24125 N$24127 N$26051 N$24246 "Waveguide Crossing" sch_x=-186 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6225 N$24129 N$24131 N$24248 N$24250 "Waveguide Crossing" sch_x=-186 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6226 N$24133 N$24135 N$24252 N$24254 "Waveguide Crossing" sch_x=-186 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6227 N$24137 N$24139 N$24256 N$24258 "Waveguide Crossing" sch_x=-186 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6228 N$24141 N$24143 N$24260 N$24262 "Waveguide Crossing" sch_x=-186 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6229 N$24145 N$24147 N$24264 N$24266 "Waveguide Crossing" sch_x=-186 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6230 N$24149 N$24151 N$24268 N$24270 "Waveguide Crossing" sch_x=-186 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6231 N$24153 N$24155 N$24272 N$24274 "Waveguide Crossing" sch_x=-186 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6232 N$24157 N$24159 N$24276 N$24278 "Waveguide Crossing" sch_x=-186 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6233 N$24161 N$24163 N$24280 N$24282 "Waveguide Crossing" sch_x=-186 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6234 N$24165 N$24167 N$24284 N$24286 "Waveguide Crossing" sch_x=-186 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6235 N$24169 N$24171 N$24288 N$24290 "Waveguide Crossing" sch_x=-186 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6236 N$24173 N$24175 N$24292 N$24294 "Waveguide Crossing" sch_x=-186 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6237 N$24177 N$24179 N$24296 N$24298 "Waveguide Crossing" sch_x=-186 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6238 N$24181 N$24183 N$24300 N$24302 "Waveguide Crossing" sch_x=-186 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6239 N$24185 N$24187 N$24304 N$24306 "Waveguide Crossing" sch_x=-186 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6240 N$24189 N$24191 N$24308 N$24310 "Waveguide Crossing" sch_x=-186 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6241 N$24193 N$24195 N$24312 N$24314 "Waveguide Crossing" sch_x=-186 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6242 N$24197 N$24199 N$24316 N$24318 "Waveguide Crossing" sch_x=-186 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6243 N$24201 N$24203 N$24320 N$24322 "Waveguide Crossing" sch_x=-186 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6244 N$24205 N$24207 N$24324 N$24326 "Waveguide Crossing" sch_x=-186 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6245 N$24209 N$24211 N$24328 N$24330 "Waveguide Crossing" sch_x=-186 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6246 N$24213 N$24215 N$24332 N$24334 "Waveguide Crossing" sch_x=-186 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6247 N$24217 N$24219 N$24336 N$24338 "Waveguide Crossing" sch_x=-186 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6248 N$24221 N$24223 N$24340 N$24342 "Waveguide Crossing" sch_x=-186 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6249 N$24225 N$24227 N$24344 N$24346 "Waveguide Crossing" sch_x=-186 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6250 N$24229 N$24231 N$24348 N$24350 "Waveguide Crossing" sch_x=-186 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6251 N$24233 N$24235 N$24352 N$24354 "Waveguide Crossing" sch_x=-186 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6252 N$24237 N$24239 N$24356 N$24358 "Waveguide Crossing" sch_x=-186 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6253 N$24241 N$24243 N$24360 N$26169 "Waveguide Crossing" sch_x=-186 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6254 N$24245 N$24247 N$26053 N$24362 "Waveguide Crossing" sch_x=-184 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6255 N$24249 N$24251 N$24364 N$24366 "Waveguide Crossing" sch_x=-184 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6256 N$24253 N$24255 N$24368 N$24370 "Waveguide Crossing" sch_x=-184 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6257 N$24257 N$24259 N$24372 N$24374 "Waveguide Crossing" sch_x=-184 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6258 N$24261 N$24263 N$24376 N$24378 "Waveguide Crossing" sch_x=-184 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6259 N$24265 N$24267 N$24380 N$24382 "Waveguide Crossing" sch_x=-184 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6260 N$24269 N$24271 N$24384 N$24386 "Waveguide Crossing" sch_x=-184 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6261 N$24273 N$24275 N$24388 N$24390 "Waveguide Crossing" sch_x=-184 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6262 N$24277 N$24279 N$24392 N$24394 "Waveguide Crossing" sch_x=-184 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6263 N$24281 N$24283 N$24396 N$24398 "Waveguide Crossing" sch_x=-184 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6264 N$24285 N$24287 N$24400 N$24402 "Waveguide Crossing" sch_x=-184 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6265 N$24289 N$24291 N$24404 N$24406 "Waveguide Crossing" sch_x=-184 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6266 N$24293 N$24295 N$24408 N$24410 "Waveguide Crossing" sch_x=-184 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6267 N$24297 N$24299 N$24412 N$24414 "Waveguide Crossing" sch_x=-184 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6268 N$24301 N$24303 N$24416 N$24418 "Waveguide Crossing" sch_x=-184 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6269 N$24305 N$24307 N$24420 N$24422 "Waveguide Crossing" sch_x=-184 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6270 N$24309 N$24311 N$24424 N$24426 "Waveguide Crossing" sch_x=-184 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6271 N$24313 N$24315 N$24428 N$24430 "Waveguide Crossing" sch_x=-184 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6272 N$24317 N$24319 N$24432 N$24434 "Waveguide Crossing" sch_x=-184 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6273 N$24321 N$24323 N$24436 N$24438 "Waveguide Crossing" sch_x=-184 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6274 N$24325 N$24327 N$24440 N$24442 "Waveguide Crossing" sch_x=-184 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6275 N$24329 N$24331 N$24444 N$24446 "Waveguide Crossing" sch_x=-184 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6276 N$24333 N$24335 N$24448 N$24450 "Waveguide Crossing" sch_x=-184 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6277 N$24337 N$24339 N$24452 N$24454 "Waveguide Crossing" sch_x=-184 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6278 N$24341 N$24343 N$24456 N$24458 "Waveguide Crossing" sch_x=-184 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6279 N$24345 N$24347 N$24460 N$24462 "Waveguide Crossing" sch_x=-184 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6280 N$24349 N$24351 N$24464 N$24466 "Waveguide Crossing" sch_x=-184 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6281 N$24353 N$24355 N$24468 N$24470 "Waveguide Crossing" sch_x=-184 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6282 N$24357 N$24359 N$24472 N$26167 "Waveguide Crossing" sch_x=-184 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6283 N$24361 N$24363 N$26055 N$24474 "Waveguide Crossing" sch_x=-182 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6284 N$24365 N$24367 N$24476 N$24478 "Waveguide Crossing" sch_x=-182 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6285 N$24369 N$24371 N$24480 N$24482 "Waveguide Crossing" sch_x=-182 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6286 N$24373 N$24375 N$24484 N$24486 "Waveguide Crossing" sch_x=-182 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6287 N$24377 N$24379 N$24488 N$24490 "Waveguide Crossing" sch_x=-182 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6288 N$24381 N$24383 N$24492 N$24494 "Waveguide Crossing" sch_x=-182 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6289 N$24385 N$24387 N$24496 N$24498 "Waveguide Crossing" sch_x=-182 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6290 N$24389 N$24391 N$24500 N$24502 "Waveguide Crossing" sch_x=-182 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6291 N$24393 N$24395 N$24504 N$24506 "Waveguide Crossing" sch_x=-182 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6292 N$24397 N$24399 N$24508 N$24510 "Waveguide Crossing" sch_x=-182 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6293 N$24401 N$24403 N$24512 N$24514 "Waveguide Crossing" sch_x=-182 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6294 N$24405 N$24407 N$24516 N$24518 "Waveguide Crossing" sch_x=-182 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6295 N$24409 N$24411 N$24520 N$24522 "Waveguide Crossing" sch_x=-182 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6296 N$24413 N$24415 N$24524 N$24526 "Waveguide Crossing" sch_x=-182 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6297 N$24417 N$24419 N$24528 N$24530 "Waveguide Crossing" sch_x=-182 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6298 N$24421 N$24423 N$24532 N$24534 "Waveguide Crossing" sch_x=-182 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6299 N$24425 N$24427 N$24536 N$24538 "Waveguide Crossing" sch_x=-182 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6300 N$24429 N$24431 N$24540 N$24542 "Waveguide Crossing" sch_x=-182 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6301 N$24433 N$24435 N$24544 N$24546 "Waveguide Crossing" sch_x=-182 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6302 N$24437 N$24439 N$24548 N$24550 "Waveguide Crossing" sch_x=-182 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6303 N$24441 N$24443 N$24552 N$24554 "Waveguide Crossing" sch_x=-182 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6304 N$24445 N$24447 N$24556 N$24558 "Waveguide Crossing" sch_x=-182 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6305 N$24449 N$24451 N$24560 N$24562 "Waveguide Crossing" sch_x=-182 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6306 N$24453 N$24455 N$24564 N$24566 "Waveguide Crossing" sch_x=-182 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6307 N$24457 N$24459 N$24568 N$24570 "Waveguide Crossing" sch_x=-182 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6308 N$24461 N$24463 N$24572 N$24574 "Waveguide Crossing" sch_x=-182 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6309 N$24465 N$24467 N$24576 N$24578 "Waveguide Crossing" sch_x=-182 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6310 N$24469 N$24471 N$24580 N$26165 "Waveguide Crossing" sch_x=-182 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6311 N$24473 N$24475 N$26057 N$24582 "Waveguide Crossing" sch_x=-180 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6312 N$24477 N$24479 N$24584 N$24586 "Waveguide Crossing" sch_x=-180 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6313 N$24481 N$24483 N$24588 N$24590 "Waveguide Crossing" sch_x=-180 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6314 N$24485 N$24487 N$24592 N$24594 "Waveguide Crossing" sch_x=-180 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6315 N$24489 N$24491 N$24596 N$24598 "Waveguide Crossing" sch_x=-180 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6316 N$24493 N$24495 N$24600 N$24602 "Waveguide Crossing" sch_x=-180 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6317 N$24497 N$24499 N$24604 N$24606 "Waveguide Crossing" sch_x=-180 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6318 N$24501 N$24503 N$24608 N$24610 "Waveguide Crossing" sch_x=-180 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6319 N$24505 N$24507 N$24612 N$24614 "Waveguide Crossing" sch_x=-180 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6320 N$24509 N$24511 N$24616 N$24618 "Waveguide Crossing" sch_x=-180 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6321 N$24513 N$24515 N$24620 N$24622 "Waveguide Crossing" sch_x=-180 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6322 N$24517 N$24519 N$24624 N$24626 "Waveguide Crossing" sch_x=-180 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6323 N$24521 N$24523 N$24628 N$24630 "Waveguide Crossing" sch_x=-180 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6324 N$24525 N$24527 N$24632 N$24634 "Waveguide Crossing" sch_x=-180 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6325 N$24529 N$24531 N$24636 N$24638 "Waveguide Crossing" sch_x=-180 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6326 N$24533 N$24535 N$24640 N$24642 "Waveguide Crossing" sch_x=-180 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6327 N$24537 N$24539 N$24644 N$24646 "Waveguide Crossing" sch_x=-180 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6328 N$24541 N$24543 N$24648 N$24650 "Waveguide Crossing" sch_x=-180 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6329 N$24545 N$24547 N$24652 N$24654 "Waveguide Crossing" sch_x=-180 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6330 N$24549 N$24551 N$24656 N$24658 "Waveguide Crossing" sch_x=-180 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6331 N$24553 N$24555 N$24660 N$24662 "Waveguide Crossing" sch_x=-180 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6332 N$24557 N$24559 N$24664 N$24666 "Waveguide Crossing" sch_x=-180 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6333 N$24561 N$24563 N$24668 N$24670 "Waveguide Crossing" sch_x=-180 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6334 N$24565 N$24567 N$24672 N$24674 "Waveguide Crossing" sch_x=-180 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6335 N$24569 N$24571 N$24676 N$24678 "Waveguide Crossing" sch_x=-180 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6336 N$24573 N$24575 N$24680 N$24682 "Waveguide Crossing" sch_x=-180 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6337 N$24577 N$24579 N$24684 N$26163 "Waveguide Crossing" sch_x=-180 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6338 N$24581 N$24583 N$26059 N$24686 "Waveguide Crossing" sch_x=-178 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6339 N$24585 N$24587 N$24688 N$24690 "Waveguide Crossing" sch_x=-178 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6340 N$24589 N$24591 N$24692 N$24694 "Waveguide Crossing" sch_x=-178 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6341 N$24593 N$24595 N$24696 N$24698 "Waveguide Crossing" sch_x=-178 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6342 N$24597 N$24599 N$24700 N$24702 "Waveguide Crossing" sch_x=-178 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6343 N$24601 N$24603 N$24704 N$24706 "Waveguide Crossing" sch_x=-178 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6344 N$24605 N$24607 N$24708 N$24710 "Waveguide Crossing" sch_x=-178 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6345 N$24609 N$24611 N$24712 N$24714 "Waveguide Crossing" sch_x=-178 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6346 N$24613 N$24615 N$24716 N$24718 "Waveguide Crossing" sch_x=-178 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6347 N$24617 N$24619 N$24720 N$24722 "Waveguide Crossing" sch_x=-178 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6348 N$24621 N$24623 N$24724 N$24726 "Waveguide Crossing" sch_x=-178 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6349 N$24625 N$24627 N$24728 N$24730 "Waveguide Crossing" sch_x=-178 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6350 N$24629 N$24631 N$24732 N$24734 "Waveguide Crossing" sch_x=-178 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6351 N$24633 N$24635 N$24736 N$24738 "Waveguide Crossing" sch_x=-178 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6352 N$24637 N$24639 N$24740 N$24742 "Waveguide Crossing" sch_x=-178 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6353 N$24641 N$24643 N$24744 N$24746 "Waveguide Crossing" sch_x=-178 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6354 N$24645 N$24647 N$24748 N$24750 "Waveguide Crossing" sch_x=-178 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6355 N$24649 N$24651 N$24752 N$24754 "Waveguide Crossing" sch_x=-178 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6356 N$24653 N$24655 N$24756 N$24758 "Waveguide Crossing" sch_x=-178 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6357 N$24657 N$24659 N$24760 N$24762 "Waveguide Crossing" sch_x=-178 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6358 N$24661 N$24663 N$24764 N$24766 "Waveguide Crossing" sch_x=-178 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6359 N$24665 N$24667 N$24768 N$24770 "Waveguide Crossing" sch_x=-178 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6360 N$24669 N$24671 N$24772 N$24774 "Waveguide Crossing" sch_x=-178 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6361 N$24673 N$24675 N$24776 N$24778 "Waveguide Crossing" sch_x=-178 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6362 N$24677 N$24679 N$24780 N$24782 "Waveguide Crossing" sch_x=-178 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6363 N$24681 N$24683 N$24784 N$26161 "Waveguide Crossing" sch_x=-178 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6364 N$24685 N$24687 N$26061 N$24786 "Waveguide Crossing" sch_x=-176 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6365 N$24689 N$24691 N$24788 N$24790 "Waveguide Crossing" sch_x=-176 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6366 N$24693 N$24695 N$24792 N$24794 "Waveguide Crossing" sch_x=-176 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6367 N$24697 N$24699 N$24796 N$24798 "Waveguide Crossing" sch_x=-176 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6368 N$24701 N$24703 N$24800 N$24802 "Waveguide Crossing" sch_x=-176 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6369 N$24705 N$24707 N$24804 N$24806 "Waveguide Crossing" sch_x=-176 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6370 N$24709 N$24711 N$24808 N$24810 "Waveguide Crossing" sch_x=-176 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6371 N$24713 N$24715 N$24812 N$24814 "Waveguide Crossing" sch_x=-176 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6372 N$24717 N$24719 N$24816 N$24818 "Waveguide Crossing" sch_x=-176 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6373 N$24721 N$24723 N$24820 N$24822 "Waveguide Crossing" sch_x=-176 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6374 N$24725 N$24727 N$24824 N$24826 "Waveguide Crossing" sch_x=-176 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6375 N$24729 N$24731 N$24828 N$24830 "Waveguide Crossing" sch_x=-176 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6376 N$24733 N$24735 N$24832 N$24834 "Waveguide Crossing" sch_x=-176 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6377 N$24737 N$24739 N$24836 N$24838 "Waveguide Crossing" sch_x=-176 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6378 N$24741 N$24743 N$24840 N$24842 "Waveguide Crossing" sch_x=-176 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6379 N$24745 N$24747 N$24844 N$24846 "Waveguide Crossing" sch_x=-176 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6380 N$24749 N$24751 N$24848 N$24850 "Waveguide Crossing" sch_x=-176 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6381 N$24753 N$24755 N$24852 N$24854 "Waveguide Crossing" sch_x=-176 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6382 N$24757 N$24759 N$24856 N$24858 "Waveguide Crossing" sch_x=-176 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6383 N$24761 N$24763 N$24860 N$24862 "Waveguide Crossing" sch_x=-176 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6384 N$24765 N$24767 N$24864 N$24866 "Waveguide Crossing" sch_x=-176 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6385 N$24769 N$24771 N$24868 N$24870 "Waveguide Crossing" sch_x=-176 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6386 N$24773 N$24775 N$24872 N$24874 "Waveguide Crossing" sch_x=-176 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6387 N$24777 N$24779 N$24876 N$24878 "Waveguide Crossing" sch_x=-176 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6388 N$24781 N$24783 N$24880 N$26159 "Waveguide Crossing" sch_x=-176 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6389 N$24785 N$24787 N$26063 N$24882 "Waveguide Crossing" sch_x=-174 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6390 N$24789 N$24791 N$24884 N$24886 "Waveguide Crossing" sch_x=-174 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6391 N$24793 N$24795 N$24888 N$24890 "Waveguide Crossing" sch_x=-174 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6392 N$24797 N$24799 N$24892 N$24894 "Waveguide Crossing" sch_x=-174 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6393 N$24801 N$24803 N$24896 N$24898 "Waveguide Crossing" sch_x=-174 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6394 N$24805 N$24807 N$24900 N$24902 "Waveguide Crossing" sch_x=-174 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6395 N$24809 N$24811 N$24904 N$24906 "Waveguide Crossing" sch_x=-174 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6396 N$24813 N$24815 N$24908 N$24910 "Waveguide Crossing" sch_x=-174 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6397 N$24817 N$24819 N$24912 N$24914 "Waveguide Crossing" sch_x=-174 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6398 N$24821 N$24823 N$24916 N$24918 "Waveguide Crossing" sch_x=-174 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6399 N$24825 N$24827 N$24920 N$24922 "Waveguide Crossing" sch_x=-174 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6400 N$24829 N$24831 N$24924 N$24926 "Waveguide Crossing" sch_x=-174 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6401 N$24833 N$24835 N$24928 N$24930 "Waveguide Crossing" sch_x=-174 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6402 N$24837 N$24839 N$24932 N$24934 "Waveguide Crossing" sch_x=-174 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6403 N$24841 N$24843 N$24936 N$24938 "Waveguide Crossing" sch_x=-174 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6404 N$24845 N$24847 N$24940 N$24942 "Waveguide Crossing" sch_x=-174 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6405 N$24849 N$24851 N$24944 N$24946 "Waveguide Crossing" sch_x=-174 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6406 N$24853 N$24855 N$24948 N$24950 "Waveguide Crossing" sch_x=-174 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6407 N$24857 N$24859 N$24952 N$24954 "Waveguide Crossing" sch_x=-174 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6408 N$24861 N$24863 N$24956 N$24958 "Waveguide Crossing" sch_x=-174 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6409 N$24865 N$24867 N$24960 N$24962 "Waveguide Crossing" sch_x=-174 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6410 N$24869 N$24871 N$24964 N$24966 "Waveguide Crossing" sch_x=-174 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6411 N$24873 N$24875 N$24968 N$24970 "Waveguide Crossing" sch_x=-174 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6412 N$24877 N$24879 N$24972 N$26157 "Waveguide Crossing" sch_x=-174 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6413 N$24881 N$24883 N$26065 N$24974 "Waveguide Crossing" sch_x=-172 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6414 N$24885 N$24887 N$24976 N$24978 "Waveguide Crossing" sch_x=-172 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6415 N$24889 N$24891 N$24980 N$24982 "Waveguide Crossing" sch_x=-172 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6416 N$24893 N$24895 N$24984 N$24986 "Waveguide Crossing" sch_x=-172 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6417 N$24897 N$24899 N$24988 N$24990 "Waveguide Crossing" sch_x=-172 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6418 N$24901 N$24903 N$24992 N$24994 "Waveguide Crossing" sch_x=-172 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6419 N$24905 N$24907 N$24996 N$24998 "Waveguide Crossing" sch_x=-172 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6420 N$24909 N$24911 N$25000 N$25002 "Waveguide Crossing" sch_x=-172 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6421 N$24913 N$24915 N$25004 N$25006 "Waveguide Crossing" sch_x=-172 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6422 N$24917 N$24919 N$25008 N$25010 "Waveguide Crossing" sch_x=-172 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6423 N$24921 N$24923 N$25012 N$25014 "Waveguide Crossing" sch_x=-172 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6424 N$24925 N$24927 N$25016 N$25018 "Waveguide Crossing" sch_x=-172 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6425 N$24929 N$24931 N$25020 N$25022 "Waveguide Crossing" sch_x=-172 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6426 N$24933 N$24935 N$25024 N$25026 "Waveguide Crossing" sch_x=-172 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6427 N$24937 N$24939 N$25028 N$25030 "Waveguide Crossing" sch_x=-172 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6428 N$24941 N$24943 N$25032 N$25034 "Waveguide Crossing" sch_x=-172 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6429 N$24945 N$24947 N$25036 N$25038 "Waveguide Crossing" sch_x=-172 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6430 N$24949 N$24951 N$25040 N$25042 "Waveguide Crossing" sch_x=-172 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6431 N$24953 N$24955 N$25044 N$25046 "Waveguide Crossing" sch_x=-172 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6432 N$24957 N$24959 N$25048 N$25050 "Waveguide Crossing" sch_x=-172 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6433 N$24961 N$24963 N$25052 N$25054 "Waveguide Crossing" sch_x=-172 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6434 N$24965 N$24967 N$25056 N$25058 "Waveguide Crossing" sch_x=-172 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6435 N$24969 N$24971 N$25060 N$26155 "Waveguide Crossing" sch_x=-172 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6436 N$24973 N$24975 N$26067 N$25062 "Waveguide Crossing" sch_x=-170 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6437 N$24977 N$24979 N$25064 N$25066 "Waveguide Crossing" sch_x=-170 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6438 N$24981 N$24983 N$25068 N$25070 "Waveguide Crossing" sch_x=-170 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6439 N$24985 N$24987 N$25072 N$25074 "Waveguide Crossing" sch_x=-170 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6440 N$24989 N$24991 N$25076 N$25078 "Waveguide Crossing" sch_x=-170 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6441 N$24993 N$24995 N$25080 N$25082 "Waveguide Crossing" sch_x=-170 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6442 N$24997 N$24999 N$25084 N$25086 "Waveguide Crossing" sch_x=-170 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6443 N$25001 N$25003 N$25088 N$25090 "Waveguide Crossing" sch_x=-170 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6444 N$25005 N$25007 N$25092 N$25094 "Waveguide Crossing" sch_x=-170 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6445 N$25009 N$25011 N$25096 N$25098 "Waveguide Crossing" sch_x=-170 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6446 N$25013 N$25015 N$25100 N$25102 "Waveguide Crossing" sch_x=-170 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6447 N$25017 N$25019 N$25104 N$25106 "Waveguide Crossing" sch_x=-170 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6448 N$25021 N$25023 N$25108 N$25110 "Waveguide Crossing" sch_x=-170 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6449 N$25025 N$25027 N$25112 N$25114 "Waveguide Crossing" sch_x=-170 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6450 N$25029 N$25031 N$25116 N$25118 "Waveguide Crossing" sch_x=-170 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6451 N$25033 N$25035 N$25120 N$25122 "Waveguide Crossing" sch_x=-170 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6452 N$25037 N$25039 N$25124 N$25126 "Waveguide Crossing" sch_x=-170 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6453 N$25041 N$25043 N$25128 N$25130 "Waveguide Crossing" sch_x=-170 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6454 N$25045 N$25047 N$25132 N$25134 "Waveguide Crossing" sch_x=-170 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6455 N$25049 N$25051 N$25136 N$25138 "Waveguide Crossing" sch_x=-170 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6456 N$25053 N$25055 N$25140 N$25142 "Waveguide Crossing" sch_x=-170 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6457 N$25057 N$25059 N$25144 N$26153 "Waveguide Crossing" sch_x=-170 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6458 N$25061 N$25063 N$26069 N$25146 "Waveguide Crossing" sch_x=-168 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6459 N$25065 N$25067 N$25148 N$25150 "Waveguide Crossing" sch_x=-168 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6460 N$25069 N$25071 N$25152 N$25154 "Waveguide Crossing" sch_x=-168 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6461 N$25073 N$25075 N$25156 N$25158 "Waveguide Crossing" sch_x=-168 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6462 N$25077 N$25079 N$25160 N$25162 "Waveguide Crossing" sch_x=-168 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6463 N$25081 N$25083 N$25164 N$25166 "Waveguide Crossing" sch_x=-168 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6464 N$25085 N$25087 N$25168 N$25170 "Waveguide Crossing" sch_x=-168 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6465 N$25089 N$25091 N$25172 N$25174 "Waveguide Crossing" sch_x=-168 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6466 N$25093 N$25095 N$25176 N$25178 "Waveguide Crossing" sch_x=-168 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6467 N$25097 N$25099 N$25180 N$25182 "Waveguide Crossing" sch_x=-168 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6468 N$25101 N$25103 N$25184 N$25186 "Waveguide Crossing" sch_x=-168 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6469 N$25105 N$25107 N$25188 N$25190 "Waveguide Crossing" sch_x=-168 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6470 N$25109 N$25111 N$25192 N$25194 "Waveguide Crossing" sch_x=-168 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6471 N$25113 N$25115 N$25196 N$25198 "Waveguide Crossing" sch_x=-168 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6472 N$25117 N$25119 N$25200 N$25202 "Waveguide Crossing" sch_x=-168 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6473 N$25121 N$25123 N$25204 N$25206 "Waveguide Crossing" sch_x=-168 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6474 N$25125 N$25127 N$25208 N$25210 "Waveguide Crossing" sch_x=-168 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6475 N$25129 N$25131 N$25212 N$25214 "Waveguide Crossing" sch_x=-168 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6476 N$25133 N$25135 N$25216 N$25218 "Waveguide Crossing" sch_x=-168 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6477 N$25137 N$25139 N$25220 N$25222 "Waveguide Crossing" sch_x=-168 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6478 N$25141 N$25143 N$25224 N$26151 "Waveguide Crossing" sch_x=-168 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6479 N$25145 N$25147 N$26071 N$25226 "Waveguide Crossing" sch_x=-166 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6480 N$25149 N$25151 N$25228 N$25230 "Waveguide Crossing" sch_x=-166 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6481 N$25153 N$25155 N$25232 N$25234 "Waveguide Crossing" sch_x=-166 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6482 N$25157 N$25159 N$25236 N$25238 "Waveguide Crossing" sch_x=-166 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6483 N$25161 N$25163 N$25240 N$25242 "Waveguide Crossing" sch_x=-166 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6484 N$25165 N$25167 N$25244 N$25246 "Waveguide Crossing" sch_x=-166 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6485 N$25169 N$25171 N$25248 N$25250 "Waveguide Crossing" sch_x=-166 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6486 N$25173 N$25175 N$25252 N$25254 "Waveguide Crossing" sch_x=-166 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6487 N$25177 N$25179 N$25256 N$25258 "Waveguide Crossing" sch_x=-166 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6488 N$25181 N$25183 N$25260 N$25262 "Waveguide Crossing" sch_x=-166 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6489 N$25185 N$25187 N$25264 N$25266 "Waveguide Crossing" sch_x=-166 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6490 N$25189 N$25191 N$25268 N$25270 "Waveguide Crossing" sch_x=-166 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6491 N$25193 N$25195 N$25272 N$25274 "Waveguide Crossing" sch_x=-166 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6492 N$25197 N$25199 N$25276 N$25278 "Waveguide Crossing" sch_x=-166 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6493 N$25201 N$25203 N$25280 N$25282 "Waveguide Crossing" sch_x=-166 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6494 N$25205 N$25207 N$25284 N$25286 "Waveguide Crossing" sch_x=-166 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6495 N$25209 N$25211 N$25288 N$25290 "Waveguide Crossing" sch_x=-166 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6496 N$25213 N$25215 N$25292 N$25294 "Waveguide Crossing" sch_x=-166 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6497 N$25217 N$25219 N$25296 N$25298 "Waveguide Crossing" sch_x=-166 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6498 N$25221 N$25223 N$25300 N$26149 "Waveguide Crossing" sch_x=-166 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6499 N$25225 N$25227 N$26073 N$25302 "Waveguide Crossing" sch_x=-164 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6500 N$25229 N$25231 N$25304 N$25306 "Waveguide Crossing" sch_x=-164 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6501 N$25233 N$25235 N$25308 N$25310 "Waveguide Crossing" sch_x=-164 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6502 N$25237 N$25239 N$25312 N$25314 "Waveguide Crossing" sch_x=-164 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6503 N$25241 N$25243 N$25316 N$25318 "Waveguide Crossing" sch_x=-164 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6504 N$25245 N$25247 N$25320 N$25322 "Waveguide Crossing" sch_x=-164 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6505 N$25249 N$25251 N$25324 N$25326 "Waveguide Crossing" sch_x=-164 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6506 N$25253 N$25255 N$25328 N$25330 "Waveguide Crossing" sch_x=-164 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6507 N$25257 N$25259 N$25332 N$25334 "Waveguide Crossing" sch_x=-164 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6508 N$25261 N$25263 N$25336 N$25338 "Waveguide Crossing" sch_x=-164 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6509 N$25265 N$25267 N$25340 N$25342 "Waveguide Crossing" sch_x=-164 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6510 N$25269 N$25271 N$25344 N$25346 "Waveguide Crossing" sch_x=-164 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6511 N$25273 N$25275 N$25348 N$25350 "Waveguide Crossing" sch_x=-164 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6512 N$25277 N$25279 N$25352 N$25354 "Waveguide Crossing" sch_x=-164 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6513 N$25281 N$25283 N$25356 N$25358 "Waveguide Crossing" sch_x=-164 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6514 N$25285 N$25287 N$25360 N$25362 "Waveguide Crossing" sch_x=-164 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6515 N$25289 N$25291 N$25364 N$25366 "Waveguide Crossing" sch_x=-164 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6516 N$25293 N$25295 N$25368 N$25370 "Waveguide Crossing" sch_x=-164 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6517 N$25297 N$25299 N$25372 N$26147 "Waveguide Crossing" sch_x=-164 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6518 N$25301 N$25303 N$26075 N$25374 "Waveguide Crossing" sch_x=-162 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6519 N$25305 N$25307 N$25376 N$25378 "Waveguide Crossing" sch_x=-162 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6520 N$25309 N$25311 N$25380 N$25382 "Waveguide Crossing" sch_x=-162 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6521 N$25313 N$25315 N$25384 N$25386 "Waveguide Crossing" sch_x=-162 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6522 N$25317 N$25319 N$25388 N$25390 "Waveguide Crossing" sch_x=-162 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6523 N$25321 N$25323 N$25392 N$25394 "Waveguide Crossing" sch_x=-162 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6524 N$25325 N$25327 N$25396 N$25398 "Waveguide Crossing" sch_x=-162 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6525 N$25329 N$25331 N$25400 N$25402 "Waveguide Crossing" sch_x=-162 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6526 N$25333 N$25335 N$25404 N$25406 "Waveguide Crossing" sch_x=-162 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6527 N$25337 N$25339 N$25408 N$25410 "Waveguide Crossing" sch_x=-162 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6528 N$25341 N$25343 N$25412 N$25414 "Waveguide Crossing" sch_x=-162 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6529 N$25345 N$25347 N$25416 N$25418 "Waveguide Crossing" sch_x=-162 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6530 N$25349 N$25351 N$25420 N$25422 "Waveguide Crossing" sch_x=-162 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6531 N$25353 N$25355 N$25424 N$25426 "Waveguide Crossing" sch_x=-162 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6532 N$25357 N$25359 N$25428 N$25430 "Waveguide Crossing" sch_x=-162 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6533 N$25361 N$25363 N$25432 N$25434 "Waveguide Crossing" sch_x=-162 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6534 N$25365 N$25367 N$25436 N$25438 "Waveguide Crossing" sch_x=-162 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6535 N$25369 N$25371 N$25440 N$26145 "Waveguide Crossing" sch_x=-162 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6536 N$25373 N$25375 N$26077 N$25442 "Waveguide Crossing" sch_x=-160 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6537 N$25377 N$25379 N$25444 N$25446 "Waveguide Crossing" sch_x=-160 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6538 N$25381 N$25383 N$25448 N$25450 "Waveguide Crossing" sch_x=-160 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6539 N$25385 N$25387 N$25452 N$25454 "Waveguide Crossing" sch_x=-160 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6540 N$25389 N$25391 N$25456 N$25458 "Waveguide Crossing" sch_x=-160 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6541 N$25393 N$25395 N$25460 N$25462 "Waveguide Crossing" sch_x=-160 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6542 N$25397 N$25399 N$25464 N$25466 "Waveguide Crossing" sch_x=-160 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6543 N$25401 N$25403 N$25468 N$25470 "Waveguide Crossing" sch_x=-160 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6544 N$25405 N$25407 N$25472 N$25474 "Waveguide Crossing" sch_x=-160 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6545 N$25409 N$25411 N$25476 N$25478 "Waveguide Crossing" sch_x=-160 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6546 N$25413 N$25415 N$25480 N$25482 "Waveguide Crossing" sch_x=-160 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6547 N$25417 N$25419 N$25484 N$25486 "Waveguide Crossing" sch_x=-160 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6548 N$25421 N$25423 N$25488 N$25490 "Waveguide Crossing" sch_x=-160 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6549 N$25425 N$25427 N$25492 N$25494 "Waveguide Crossing" sch_x=-160 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6550 N$25429 N$25431 N$25496 N$25498 "Waveguide Crossing" sch_x=-160 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6551 N$25433 N$25435 N$25500 N$25502 "Waveguide Crossing" sch_x=-160 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6552 N$25437 N$25439 N$25504 N$26143 "Waveguide Crossing" sch_x=-160 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6553 N$25441 N$25443 N$26079 N$25506 "Waveguide Crossing" sch_x=-158 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6554 N$25445 N$25447 N$25508 N$25510 "Waveguide Crossing" sch_x=-158 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6555 N$25449 N$25451 N$25512 N$25514 "Waveguide Crossing" sch_x=-158 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6556 N$25453 N$25455 N$25516 N$25518 "Waveguide Crossing" sch_x=-158 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6557 N$25457 N$25459 N$25520 N$25522 "Waveguide Crossing" sch_x=-158 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6558 N$25461 N$25463 N$25524 N$25526 "Waveguide Crossing" sch_x=-158 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6559 N$25465 N$25467 N$25528 N$25530 "Waveguide Crossing" sch_x=-158 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6560 N$25469 N$25471 N$25532 N$25534 "Waveguide Crossing" sch_x=-158 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6561 N$25473 N$25475 N$25536 N$25538 "Waveguide Crossing" sch_x=-158 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6562 N$25477 N$25479 N$25540 N$25542 "Waveguide Crossing" sch_x=-158 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6563 N$25481 N$25483 N$25544 N$25546 "Waveguide Crossing" sch_x=-158 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6564 N$25485 N$25487 N$25548 N$25550 "Waveguide Crossing" sch_x=-158 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6565 N$25489 N$25491 N$25552 N$25554 "Waveguide Crossing" sch_x=-158 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6566 N$25493 N$25495 N$25556 N$25558 "Waveguide Crossing" sch_x=-158 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6567 N$25497 N$25499 N$25560 N$25562 "Waveguide Crossing" sch_x=-158 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6568 N$25501 N$25503 N$25564 N$26141 "Waveguide Crossing" sch_x=-158 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6569 N$25505 N$25507 N$26081 N$25566 "Waveguide Crossing" sch_x=-156 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6570 N$25509 N$25511 N$25568 N$25570 "Waveguide Crossing" sch_x=-156 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6571 N$25513 N$25515 N$25572 N$25574 "Waveguide Crossing" sch_x=-156 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6572 N$25517 N$25519 N$25576 N$25578 "Waveguide Crossing" sch_x=-156 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6573 N$25521 N$25523 N$25580 N$25582 "Waveguide Crossing" sch_x=-156 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6574 N$25525 N$25527 N$25584 N$25586 "Waveguide Crossing" sch_x=-156 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6575 N$25529 N$25531 N$25588 N$25590 "Waveguide Crossing" sch_x=-156 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6576 N$25533 N$25535 N$25592 N$25594 "Waveguide Crossing" sch_x=-156 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6577 N$25537 N$25539 N$25596 N$25598 "Waveguide Crossing" sch_x=-156 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6578 N$25541 N$25543 N$25600 N$25602 "Waveguide Crossing" sch_x=-156 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6579 N$25545 N$25547 N$25604 N$25606 "Waveguide Crossing" sch_x=-156 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6580 N$25549 N$25551 N$25608 N$25610 "Waveguide Crossing" sch_x=-156 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6581 N$25553 N$25555 N$25612 N$25614 "Waveguide Crossing" sch_x=-156 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6582 N$25557 N$25559 N$25616 N$25618 "Waveguide Crossing" sch_x=-156 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6583 N$25561 N$25563 N$25620 N$26139 "Waveguide Crossing" sch_x=-156 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6584 N$25565 N$25567 N$26083 N$25622 "Waveguide Crossing" sch_x=-154 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6585 N$25569 N$25571 N$25624 N$25626 "Waveguide Crossing" sch_x=-154 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6586 N$25573 N$25575 N$25628 N$25630 "Waveguide Crossing" sch_x=-154 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6587 N$25577 N$25579 N$25632 N$25634 "Waveguide Crossing" sch_x=-154 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6588 N$25581 N$25583 N$25636 N$25638 "Waveguide Crossing" sch_x=-154 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6589 N$25585 N$25587 N$25640 N$25642 "Waveguide Crossing" sch_x=-154 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6590 N$25589 N$25591 N$25644 N$25646 "Waveguide Crossing" sch_x=-154 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6591 N$25593 N$25595 N$25648 N$25650 "Waveguide Crossing" sch_x=-154 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6592 N$25597 N$25599 N$25652 N$25654 "Waveguide Crossing" sch_x=-154 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6593 N$25601 N$25603 N$25656 N$25658 "Waveguide Crossing" sch_x=-154 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6594 N$25605 N$25607 N$25660 N$25662 "Waveguide Crossing" sch_x=-154 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6595 N$25609 N$25611 N$25664 N$25666 "Waveguide Crossing" sch_x=-154 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6596 N$25613 N$25615 N$25668 N$25670 "Waveguide Crossing" sch_x=-154 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6597 N$25617 N$25619 N$25672 N$26137 "Waveguide Crossing" sch_x=-154 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6598 N$25621 N$25623 N$26085 N$25674 "Waveguide Crossing" sch_x=-152 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6599 N$25625 N$25627 N$25676 N$25678 "Waveguide Crossing" sch_x=-152 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6600 N$25629 N$25631 N$25680 N$25682 "Waveguide Crossing" sch_x=-152 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6601 N$25633 N$25635 N$25684 N$25686 "Waveguide Crossing" sch_x=-152 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6602 N$25637 N$25639 N$25688 N$25690 "Waveguide Crossing" sch_x=-152 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6603 N$25641 N$25643 N$25692 N$25694 "Waveguide Crossing" sch_x=-152 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6604 N$25645 N$25647 N$25696 N$25698 "Waveguide Crossing" sch_x=-152 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6605 N$25649 N$25651 N$25700 N$25702 "Waveguide Crossing" sch_x=-152 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6606 N$25653 N$25655 N$25704 N$25706 "Waveguide Crossing" sch_x=-152 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6607 N$25657 N$25659 N$25708 N$25710 "Waveguide Crossing" sch_x=-152 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6608 N$25661 N$25663 N$25712 N$25714 "Waveguide Crossing" sch_x=-152 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6609 N$25665 N$25667 N$25716 N$25718 "Waveguide Crossing" sch_x=-152 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6610 N$25669 N$25671 N$25720 N$26135 "Waveguide Crossing" sch_x=-152 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6611 N$25673 N$25675 N$26087 N$25722 "Waveguide Crossing" sch_x=-150 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6612 N$25677 N$25679 N$25724 N$25726 "Waveguide Crossing" sch_x=-150 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6613 N$25681 N$25683 N$25728 N$25730 "Waveguide Crossing" sch_x=-150 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6614 N$25685 N$25687 N$25732 N$25734 "Waveguide Crossing" sch_x=-150 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6615 N$25689 N$25691 N$25736 N$25738 "Waveguide Crossing" sch_x=-150 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6616 N$25693 N$25695 N$25740 N$25742 "Waveguide Crossing" sch_x=-150 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6617 N$25697 N$25699 N$25744 N$25746 "Waveguide Crossing" sch_x=-150 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6618 N$25701 N$25703 N$25748 N$25750 "Waveguide Crossing" sch_x=-150 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6619 N$25705 N$25707 N$25752 N$25754 "Waveguide Crossing" sch_x=-150 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6620 N$25709 N$25711 N$25756 N$25758 "Waveguide Crossing" sch_x=-150 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6621 N$25713 N$25715 N$25760 N$25762 "Waveguide Crossing" sch_x=-150 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6622 N$25717 N$25719 N$25764 N$26133 "Waveguide Crossing" sch_x=-150 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6623 N$25721 N$25723 N$26089 N$25766 "Waveguide Crossing" sch_x=-148 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6624 N$25725 N$25727 N$25768 N$25770 "Waveguide Crossing" sch_x=-148 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6625 N$25729 N$25731 N$25772 N$25774 "Waveguide Crossing" sch_x=-148 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6626 N$25733 N$25735 N$25776 N$25778 "Waveguide Crossing" sch_x=-148 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6627 N$25737 N$25739 N$25780 N$25782 "Waveguide Crossing" sch_x=-148 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6628 N$25741 N$25743 N$25784 N$25786 "Waveguide Crossing" sch_x=-148 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6629 N$25745 N$25747 N$25788 N$25790 "Waveguide Crossing" sch_x=-148 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6630 N$25749 N$25751 N$25792 N$25794 "Waveguide Crossing" sch_x=-148 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6631 N$25753 N$25755 N$25796 N$25798 "Waveguide Crossing" sch_x=-148 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6632 N$25757 N$25759 N$25800 N$25802 "Waveguide Crossing" sch_x=-148 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6633 N$25761 N$25763 N$25804 N$26131 "Waveguide Crossing" sch_x=-148 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6634 N$25765 N$25767 N$26091 N$25806 "Waveguide Crossing" sch_x=-146 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6635 N$25769 N$25771 N$25808 N$25810 "Waveguide Crossing" sch_x=-146 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6636 N$25773 N$25775 N$25812 N$25814 "Waveguide Crossing" sch_x=-146 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6637 N$25777 N$25779 N$25816 N$25818 "Waveguide Crossing" sch_x=-146 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6638 N$25781 N$25783 N$25820 N$25822 "Waveguide Crossing" sch_x=-146 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6639 N$25785 N$25787 N$25824 N$25826 "Waveguide Crossing" sch_x=-146 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6640 N$25789 N$25791 N$25828 N$25830 "Waveguide Crossing" sch_x=-146 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6641 N$25793 N$25795 N$25832 N$25834 "Waveguide Crossing" sch_x=-146 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6642 N$25797 N$25799 N$25836 N$25838 "Waveguide Crossing" sch_x=-146 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6643 N$25801 N$25803 N$25840 N$26129 "Waveguide Crossing" sch_x=-146 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6644 N$25805 N$25807 N$26093 N$25842 "Waveguide Crossing" sch_x=-144 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6645 N$25809 N$25811 N$25844 N$25846 "Waveguide Crossing" sch_x=-144 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6646 N$25813 N$25815 N$25848 N$25850 "Waveguide Crossing" sch_x=-144 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6647 N$25817 N$25819 N$25852 N$25854 "Waveguide Crossing" sch_x=-144 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6648 N$25821 N$25823 N$25856 N$25858 "Waveguide Crossing" sch_x=-144 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6649 N$25825 N$25827 N$25860 N$25862 "Waveguide Crossing" sch_x=-144 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6650 N$25829 N$25831 N$25864 N$25866 "Waveguide Crossing" sch_x=-144 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6651 N$25833 N$25835 N$25868 N$25870 "Waveguide Crossing" sch_x=-144 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6652 N$25837 N$25839 N$25872 N$26127 "Waveguide Crossing" sch_x=-144 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6653 N$25841 N$25843 N$26095 N$25874 "Waveguide Crossing" sch_x=-142 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6654 N$25845 N$25847 N$25876 N$25878 "Waveguide Crossing" sch_x=-142 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6655 N$25849 N$25851 N$25880 N$25882 "Waveguide Crossing" sch_x=-142 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6656 N$25853 N$25855 N$25884 N$25886 "Waveguide Crossing" sch_x=-142 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6657 N$25857 N$25859 N$25888 N$25890 "Waveguide Crossing" sch_x=-142 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6658 N$25861 N$25863 N$25892 N$25894 "Waveguide Crossing" sch_x=-142 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6659 N$25865 N$25867 N$25896 N$25898 "Waveguide Crossing" sch_x=-142 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6660 N$25869 N$25871 N$25900 N$26125 "Waveguide Crossing" sch_x=-142 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6661 N$25873 N$25875 N$26097 N$25902 "Waveguide Crossing" sch_x=-140 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6662 N$25877 N$25879 N$25904 N$25906 "Waveguide Crossing" sch_x=-140 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6663 N$25881 N$25883 N$25908 N$25910 "Waveguide Crossing" sch_x=-140 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6664 N$25885 N$25887 N$25912 N$25914 "Waveguide Crossing" sch_x=-140 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6665 N$25889 N$25891 N$25916 N$25918 "Waveguide Crossing" sch_x=-140 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6666 N$25893 N$25895 N$25920 N$25922 "Waveguide Crossing" sch_x=-140 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6667 N$25897 N$25899 N$25924 N$26123 "Waveguide Crossing" sch_x=-140 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6668 N$25901 N$25903 N$26099 N$25926 "Waveguide Crossing" sch_x=-138 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6669 N$25905 N$25907 N$25928 N$25930 "Waveguide Crossing" sch_x=-138 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6670 N$25909 N$25911 N$25932 N$25934 "Waveguide Crossing" sch_x=-138 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6671 N$25913 N$25915 N$25936 N$25938 "Waveguide Crossing" sch_x=-138 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6672 N$25917 N$25919 N$25940 N$25942 "Waveguide Crossing" sch_x=-138 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6673 N$25921 N$25923 N$25944 N$26121 "Waveguide Crossing" sch_x=-138 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6674 N$25925 N$25927 N$26101 N$25946 "Waveguide Crossing" sch_x=-136 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6675 N$25929 N$25931 N$25948 N$25950 "Waveguide Crossing" sch_x=-136 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6676 N$25933 N$25935 N$25952 N$25954 "Waveguide Crossing" sch_x=-136 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6677 N$25937 N$25939 N$25956 N$25958 "Waveguide Crossing" sch_x=-136 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6678 N$25941 N$25943 N$25960 N$26119 "Waveguide Crossing" sch_x=-136 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6679 N$25945 N$25947 N$26103 N$25962 "Waveguide Crossing" sch_x=-134 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6680 N$25949 N$25951 N$25964 N$25966 "Waveguide Crossing" sch_x=-134 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6681 N$25953 N$25955 N$25968 N$25970 "Waveguide Crossing" sch_x=-134 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6682 N$25957 N$25959 N$25972 N$26117 "Waveguide Crossing" sch_x=-134 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6683 N$25961 N$25963 N$26105 N$25974 "Waveguide Crossing" sch_x=-132 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6684 N$25965 N$25967 N$25976 N$25978 "Waveguide Crossing" sch_x=-132 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6685 N$25969 N$25971 N$25980 N$26115 "Waveguide Crossing" sch_x=-132 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6686 N$25973 N$25975 N$26107 N$25982 "Waveguide Crossing" sch_x=-130 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6687 N$25977 N$25979 N$25984 N$26113 "Waveguide Crossing" sch_x=-130 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6688 N$25981 N$25983 N$26109 N$26111 "Waveguide Crossing" sch_x=-128 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3553 N$26112 N$26114 N$15805 N$13698 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3554 N$26116 N$26118 N$13700 N$13702 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3555 N$26120 N$26122 N$13704 N$13706 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3556 N$26124 N$26126 N$13708 N$13710 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3557 N$26128 N$26130 N$13712 N$13714 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3558 N$26132 N$26134 N$13716 N$13718 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3559 N$26136 N$26138 N$13720 N$13722 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3560 N$26140 N$26142 N$13724 N$13726 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3561 N$26144 N$26146 N$13728 N$13730 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3562 N$26148 N$26150 N$13732 N$13734 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3563 N$26152 N$26154 N$13736 N$13738 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3564 N$26156 N$26158 N$13740 N$13742 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3565 N$26160 N$26162 N$13744 N$13746 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3566 N$26164 N$26166 N$13748 N$13750 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3567 N$26168 N$26170 N$13752 N$13754 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3568 N$26172 N$26174 N$13756 N$13758 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3569 N$26176 N$26178 N$13760 N$13762 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3570 N$26180 N$26182 N$13764 N$13766 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3571 N$26184 N$26186 N$13768 N$13770 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3572 N$26188 N$26190 N$13772 N$13774 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3573 N$26192 N$26194 N$13776 N$13778 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3574 N$26196 N$26198 N$13780 N$13782 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3575 N$26200 N$26202 N$13784 N$13786 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3576 N$26204 N$26206 N$13788 N$13790 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3577 N$26208 N$26210 N$13792 N$13794 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3578 N$26212 N$26214 N$13796 N$13798 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3579 N$26216 N$26218 N$13800 N$13802 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3580 N$26220 N$26222 N$13804 N$13806 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3581 N$26224 N$26226 N$13808 N$13810 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3582 N$26228 N$26230 N$13812 N$13814 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3583 N$26232 N$26234 N$13816 N$13818 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3584 N$26236 N$26240 N$13820 N$15807 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3585 N$13697 N$13699 N$15681 N$13822 "Waveguide Crossing" sch_x=-124 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3586 N$13701 N$13703 N$13824 N$13826 "Waveguide Crossing" sch_x=-124 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3587 N$13705 N$13707 N$13828 N$13830 "Waveguide Crossing" sch_x=-124 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3588 N$13709 N$13711 N$13832 N$13834 "Waveguide Crossing" sch_x=-124 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3589 N$13713 N$13715 N$13836 N$13838 "Waveguide Crossing" sch_x=-124 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3590 N$13717 N$13719 N$13840 N$13842 "Waveguide Crossing" sch_x=-124 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3591 N$13721 N$13723 N$13844 N$13846 "Waveguide Crossing" sch_x=-124 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3592 N$13725 N$13727 N$13848 N$13850 "Waveguide Crossing" sch_x=-124 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3593 N$13729 N$13731 N$13852 N$13854 "Waveguide Crossing" sch_x=-124 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3594 N$13733 N$13735 N$13856 N$13858 "Waveguide Crossing" sch_x=-124 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3595 N$13737 N$13739 N$13860 N$13862 "Waveguide Crossing" sch_x=-124 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3596 N$13741 N$13743 N$13864 N$13866 "Waveguide Crossing" sch_x=-124 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3597 N$13745 N$13747 N$13868 N$13870 "Waveguide Crossing" sch_x=-124 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3598 N$13749 N$13751 N$13872 N$13874 "Waveguide Crossing" sch_x=-124 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3599 N$13753 N$13755 N$13876 N$13878 "Waveguide Crossing" sch_x=-124 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3600 N$13757 N$13759 N$13880 N$13882 "Waveguide Crossing" sch_x=-124 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3601 N$13761 N$13763 N$13884 N$13886 "Waveguide Crossing" sch_x=-124 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3602 N$13765 N$13767 N$13888 N$13890 "Waveguide Crossing" sch_x=-124 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3603 N$13769 N$13771 N$13892 N$13894 "Waveguide Crossing" sch_x=-124 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3604 N$13773 N$13775 N$13896 N$13898 "Waveguide Crossing" sch_x=-124 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3605 N$13777 N$13779 N$13900 N$13902 "Waveguide Crossing" sch_x=-124 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3606 N$13781 N$13783 N$13904 N$13906 "Waveguide Crossing" sch_x=-124 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3607 N$13785 N$13787 N$13908 N$13910 "Waveguide Crossing" sch_x=-124 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3608 N$13789 N$13791 N$13912 N$13914 "Waveguide Crossing" sch_x=-124 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3609 N$13793 N$13795 N$13916 N$13918 "Waveguide Crossing" sch_x=-124 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3610 N$13797 N$13799 N$13920 N$13922 "Waveguide Crossing" sch_x=-124 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3611 N$13801 N$13803 N$13924 N$13926 "Waveguide Crossing" sch_x=-124 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3612 N$13805 N$13807 N$13928 N$13930 "Waveguide Crossing" sch_x=-124 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3613 N$13809 N$13811 N$13932 N$13934 "Waveguide Crossing" sch_x=-124 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3614 N$13813 N$13815 N$13936 N$13938 "Waveguide Crossing" sch_x=-124 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3615 N$13817 N$13819 N$13940 N$15803 "Waveguide Crossing" sch_x=-124 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3616 N$13821 N$13823 N$15683 N$13942 "Waveguide Crossing" sch_x=-122 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3617 N$13825 N$13827 N$13944 N$13946 "Waveguide Crossing" sch_x=-122 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3618 N$13829 N$13831 N$13948 N$13950 "Waveguide Crossing" sch_x=-122 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3619 N$13833 N$13835 N$13952 N$13954 "Waveguide Crossing" sch_x=-122 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3620 N$13837 N$13839 N$13956 N$13958 "Waveguide Crossing" sch_x=-122 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3621 N$13841 N$13843 N$13960 N$13962 "Waveguide Crossing" sch_x=-122 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3622 N$13845 N$13847 N$13964 N$13966 "Waveguide Crossing" sch_x=-122 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3623 N$13849 N$13851 N$13968 N$13970 "Waveguide Crossing" sch_x=-122 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3624 N$13853 N$13855 N$13972 N$13974 "Waveguide Crossing" sch_x=-122 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3625 N$13857 N$13859 N$13976 N$13978 "Waveguide Crossing" sch_x=-122 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3626 N$13861 N$13863 N$13980 N$13982 "Waveguide Crossing" sch_x=-122 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3627 N$13865 N$13867 N$13984 N$13986 "Waveguide Crossing" sch_x=-122 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3628 N$13869 N$13871 N$13988 N$13990 "Waveguide Crossing" sch_x=-122 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3629 N$13873 N$13875 N$13992 N$13994 "Waveguide Crossing" sch_x=-122 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3630 N$13877 N$13879 N$13996 N$13998 "Waveguide Crossing" sch_x=-122 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3631 N$13881 N$13883 N$14000 N$14002 "Waveguide Crossing" sch_x=-122 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3632 N$13885 N$13887 N$14004 N$14006 "Waveguide Crossing" sch_x=-122 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3633 N$13889 N$13891 N$14008 N$14010 "Waveguide Crossing" sch_x=-122 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3634 N$13893 N$13895 N$14012 N$14014 "Waveguide Crossing" sch_x=-122 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3635 N$13897 N$13899 N$14016 N$14018 "Waveguide Crossing" sch_x=-122 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3636 N$13901 N$13903 N$14020 N$14022 "Waveguide Crossing" sch_x=-122 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3637 N$13905 N$13907 N$14024 N$14026 "Waveguide Crossing" sch_x=-122 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3638 N$13909 N$13911 N$14028 N$14030 "Waveguide Crossing" sch_x=-122 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3639 N$13913 N$13915 N$14032 N$14034 "Waveguide Crossing" sch_x=-122 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3640 N$13917 N$13919 N$14036 N$14038 "Waveguide Crossing" sch_x=-122 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3641 N$13921 N$13923 N$14040 N$14042 "Waveguide Crossing" sch_x=-122 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3642 N$13925 N$13927 N$14044 N$14046 "Waveguide Crossing" sch_x=-122 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3643 N$13929 N$13931 N$14048 N$14050 "Waveguide Crossing" sch_x=-122 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3644 N$13933 N$13935 N$14052 N$14054 "Waveguide Crossing" sch_x=-122 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3645 N$13937 N$13939 N$14056 N$15801 "Waveguide Crossing" sch_x=-122 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3646 N$13941 N$13943 N$15685 N$14058 "Waveguide Crossing" sch_x=-120 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3647 N$13945 N$13947 N$14060 N$14062 "Waveguide Crossing" sch_x=-120 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3648 N$13949 N$13951 N$14064 N$14066 "Waveguide Crossing" sch_x=-120 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3649 N$13953 N$13955 N$14068 N$14070 "Waveguide Crossing" sch_x=-120 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3650 N$13957 N$13959 N$14072 N$14074 "Waveguide Crossing" sch_x=-120 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3651 N$13961 N$13963 N$14076 N$14078 "Waveguide Crossing" sch_x=-120 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3652 N$13965 N$13967 N$14080 N$14082 "Waveguide Crossing" sch_x=-120 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3653 N$13969 N$13971 N$14084 N$14086 "Waveguide Crossing" sch_x=-120 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3654 N$13973 N$13975 N$14088 N$14090 "Waveguide Crossing" sch_x=-120 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3655 N$13977 N$13979 N$14092 N$14094 "Waveguide Crossing" sch_x=-120 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3656 N$13981 N$13983 N$14096 N$14098 "Waveguide Crossing" sch_x=-120 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3657 N$13985 N$13987 N$14100 N$14102 "Waveguide Crossing" sch_x=-120 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3658 N$13989 N$13991 N$14104 N$14106 "Waveguide Crossing" sch_x=-120 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3659 N$13993 N$13995 N$14108 N$14110 "Waveguide Crossing" sch_x=-120 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3660 N$13997 N$13999 N$14112 N$14114 "Waveguide Crossing" sch_x=-120 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3661 N$14001 N$14003 N$14116 N$14118 "Waveguide Crossing" sch_x=-120 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3662 N$14005 N$14007 N$14120 N$14122 "Waveguide Crossing" sch_x=-120 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3663 N$14009 N$14011 N$14124 N$14126 "Waveguide Crossing" sch_x=-120 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3664 N$14013 N$14015 N$14128 N$14130 "Waveguide Crossing" sch_x=-120 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3665 N$14017 N$14019 N$14132 N$14134 "Waveguide Crossing" sch_x=-120 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3666 N$14021 N$14023 N$14136 N$14138 "Waveguide Crossing" sch_x=-120 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3667 N$14025 N$14027 N$14140 N$14142 "Waveguide Crossing" sch_x=-120 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3668 N$14029 N$14031 N$14144 N$14146 "Waveguide Crossing" sch_x=-120 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3669 N$14033 N$14035 N$14148 N$14150 "Waveguide Crossing" sch_x=-120 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3670 N$14037 N$14039 N$14152 N$14154 "Waveguide Crossing" sch_x=-120 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3671 N$14041 N$14043 N$14156 N$14158 "Waveguide Crossing" sch_x=-120 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3672 N$14045 N$14047 N$14160 N$14162 "Waveguide Crossing" sch_x=-120 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3673 N$14049 N$14051 N$14164 N$14166 "Waveguide Crossing" sch_x=-120 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3674 N$14053 N$14055 N$14168 N$15799 "Waveguide Crossing" sch_x=-120 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3675 N$14057 N$14059 N$15687 N$14170 "Waveguide Crossing" sch_x=-118 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3676 N$14061 N$14063 N$14172 N$14174 "Waveguide Crossing" sch_x=-118 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3677 N$14065 N$14067 N$14176 N$14178 "Waveguide Crossing" sch_x=-118 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3678 N$14069 N$14071 N$14180 N$14182 "Waveguide Crossing" sch_x=-118 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3679 N$14073 N$14075 N$14184 N$14186 "Waveguide Crossing" sch_x=-118 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3680 N$14077 N$14079 N$14188 N$14190 "Waveguide Crossing" sch_x=-118 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3681 N$14081 N$14083 N$14192 N$14194 "Waveguide Crossing" sch_x=-118 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3682 N$14085 N$14087 N$14196 N$14198 "Waveguide Crossing" sch_x=-118 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3683 N$14089 N$14091 N$14200 N$14202 "Waveguide Crossing" sch_x=-118 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3684 N$14093 N$14095 N$14204 N$14206 "Waveguide Crossing" sch_x=-118 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3685 N$14097 N$14099 N$14208 N$14210 "Waveguide Crossing" sch_x=-118 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3686 N$14101 N$14103 N$14212 N$14214 "Waveguide Crossing" sch_x=-118 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3687 N$14105 N$14107 N$14216 N$14218 "Waveguide Crossing" sch_x=-118 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3688 N$14109 N$14111 N$14220 N$14222 "Waveguide Crossing" sch_x=-118 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3689 N$14113 N$14115 N$14224 N$14226 "Waveguide Crossing" sch_x=-118 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3690 N$14117 N$14119 N$14228 N$14230 "Waveguide Crossing" sch_x=-118 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3691 N$14121 N$14123 N$14232 N$14234 "Waveguide Crossing" sch_x=-118 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3692 N$14125 N$14127 N$14236 N$14238 "Waveguide Crossing" sch_x=-118 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3693 N$14129 N$14131 N$14240 N$14242 "Waveguide Crossing" sch_x=-118 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3694 N$14133 N$14135 N$14244 N$14246 "Waveguide Crossing" sch_x=-118 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3695 N$14137 N$14139 N$14248 N$14250 "Waveguide Crossing" sch_x=-118 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3696 N$14141 N$14143 N$14252 N$14254 "Waveguide Crossing" sch_x=-118 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3697 N$14145 N$14147 N$14256 N$14258 "Waveguide Crossing" sch_x=-118 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3698 N$14149 N$14151 N$14260 N$14262 "Waveguide Crossing" sch_x=-118 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3699 N$14153 N$14155 N$14264 N$14266 "Waveguide Crossing" sch_x=-118 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3700 N$14157 N$14159 N$14268 N$14270 "Waveguide Crossing" sch_x=-118 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3701 N$14161 N$14163 N$14272 N$14274 "Waveguide Crossing" sch_x=-118 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3702 N$14165 N$14167 N$14276 N$15797 "Waveguide Crossing" sch_x=-118 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3703 N$14169 N$14171 N$15689 N$14278 "Waveguide Crossing" sch_x=-116 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3704 N$14173 N$14175 N$14280 N$14282 "Waveguide Crossing" sch_x=-116 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3705 N$14177 N$14179 N$14284 N$14286 "Waveguide Crossing" sch_x=-116 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3706 N$14181 N$14183 N$14288 N$14290 "Waveguide Crossing" sch_x=-116 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3707 N$14185 N$14187 N$14292 N$14294 "Waveguide Crossing" sch_x=-116 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3708 N$14189 N$14191 N$14296 N$14298 "Waveguide Crossing" sch_x=-116 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3709 N$14193 N$14195 N$14300 N$14302 "Waveguide Crossing" sch_x=-116 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3710 N$14197 N$14199 N$14304 N$14306 "Waveguide Crossing" sch_x=-116 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3711 N$14201 N$14203 N$14308 N$14310 "Waveguide Crossing" sch_x=-116 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3712 N$14205 N$14207 N$14312 N$14314 "Waveguide Crossing" sch_x=-116 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3713 N$14209 N$14211 N$14316 N$14318 "Waveguide Crossing" sch_x=-116 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3714 N$14213 N$14215 N$14320 N$14322 "Waveguide Crossing" sch_x=-116 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3715 N$14217 N$14219 N$14324 N$14326 "Waveguide Crossing" sch_x=-116 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3716 N$14221 N$14223 N$14328 N$14330 "Waveguide Crossing" sch_x=-116 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3717 N$14225 N$14227 N$14332 N$14334 "Waveguide Crossing" sch_x=-116 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3718 N$14229 N$14231 N$14336 N$14338 "Waveguide Crossing" sch_x=-116 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3719 N$14233 N$14235 N$14340 N$14342 "Waveguide Crossing" sch_x=-116 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3720 N$14237 N$14239 N$14344 N$14346 "Waveguide Crossing" sch_x=-116 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3721 N$14241 N$14243 N$14348 N$14350 "Waveguide Crossing" sch_x=-116 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3722 N$14245 N$14247 N$14352 N$14354 "Waveguide Crossing" sch_x=-116 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3723 N$14249 N$14251 N$14356 N$14358 "Waveguide Crossing" sch_x=-116 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3724 N$14253 N$14255 N$14360 N$14362 "Waveguide Crossing" sch_x=-116 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3725 N$14257 N$14259 N$14364 N$14366 "Waveguide Crossing" sch_x=-116 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3726 N$14261 N$14263 N$14368 N$14370 "Waveguide Crossing" sch_x=-116 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3727 N$14265 N$14267 N$14372 N$14374 "Waveguide Crossing" sch_x=-116 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3728 N$14269 N$14271 N$14376 N$14378 "Waveguide Crossing" sch_x=-116 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3729 N$14273 N$14275 N$14380 N$15795 "Waveguide Crossing" sch_x=-116 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3730 N$14277 N$14279 N$15691 N$14382 "Waveguide Crossing" sch_x=-114 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3731 N$14281 N$14283 N$14384 N$14386 "Waveguide Crossing" sch_x=-114 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3732 N$14285 N$14287 N$14388 N$14390 "Waveguide Crossing" sch_x=-114 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3733 N$14289 N$14291 N$14392 N$14394 "Waveguide Crossing" sch_x=-114 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3734 N$14293 N$14295 N$14396 N$14398 "Waveguide Crossing" sch_x=-114 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3735 N$14297 N$14299 N$14400 N$14402 "Waveguide Crossing" sch_x=-114 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3736 N$14301 N$14303 N$14404 N$14406 "Waveguide Crossing" sch_x=-114 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3737 N$14305 N$14307 N$14408 N$14410 "Waveguide Crossing" sch_x=-114 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3738 N$14309 N$14311 N$14412 N$14414 "Waveguide Crossing" sch_x=-114 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3739 N$14313 N$14315 N$14416 N$14418 "Waveguide Crossing" sch_x=-114 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3740 N$14317 N$14319 N$14420 N$14422 "Waveguide Crossing" sch_x=-114 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3741 N$14321 N$14323 N$14424 N$14426 "Waveguide Crossing" sch_x=-114 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3742 N$14325 N$14327 N$14428 N$14430 "Waveguide Crossing" sch_x=-114 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3743 N$14329 N$14331 N$14432 N$14434 "Waveguide Crossing" sch_x=-114 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3744 N$14333 N$14335 N$14436 N$14438 "Waveguide Crossing" sch_x=-114 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3745 N$14337 N$14339 N$14440 N$14442 "Waveguide Crossing" sch_x=-114 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3746 N$14341 N$14343 N$14444 N$14446 "Waveguide Crossing" sch_x=-114 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3747 N$14345 N$14347 N$14448 N$14450 "Waveguide Crossing" sch_x=-114 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3748 N$14349 N$14351 N$14452 N$14454 "Waveguide Crossing" sch_x=-114 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3749 N$14353 N$14355 N$14456 N$14458 "Waveguide Crossing" sch_x=-114 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3750 N$14357 N$14359 N$14460 N$14462 "Waveguide Crossing" sch_x=-114 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3751 N$14361 N$14363 N$14464 N$14466 "Waveguide Crossing" sch_x=-114 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3752 N$14365 N$14367 N$14468 N$14470 "Waveguide Crossing" sch_x=-114 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3753 N$14369 N$14371 N$14472 N$14474 "Waveguide Crossing" sch_x=-114 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3754 N$14373 N$14375 N$14476 N$14478 "Waveguide Crossing" sch_x=-114 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3755 N$14377 N$14379 N$14480 N$15793 "Waveguide Crossing" sch_x=-114 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3756 N$14381 N$14383 N$15693 N$14482 "Waveguide Crossing" sch_x=-112 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3757 N$14385 N$14387 N$14484 N$14486 "Waveguide Crossing" sch_x=-112 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3758 N$14389 N$14391 N$14488 N$14490 "Waveguide Crossing" sch_x=-112 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3759 N$14393 N$14395 N$14492 N$14494 "Waveguide Crossing" sch_x=-112 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3760 N$14397 N$14399 N$14496 N$14498 "Waveguide Crossing" sch_x=-112 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3761 N$14401 N$14403 N$14500 N$14502 "Waveguide Crossing" sch_x=-112 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3762 N$14405 N$14407 N$14504 N$14506 "Waveguide Crossing" sch_x=-112 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3763 N$14409 N$14411 N$14508 N$14510 "Waveguide Crossing" sch_x=-112 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3764 N$14413 N$14415 N$14512 N$14514 "Waveguide Crossing" sch_x=-112 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3765 N$14417 N$14419 N$14516 N$14518 "Waveguide Crossing" sch_x=-112 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3766 N$14421 N$14423 N$14520 N$14522 "Waveguide Crossing" sch_x=-112 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3767 N$14425 N$14427 N$14524 N$14526 "Waveguide Crossing" sch_x=-112 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3768 N$14429 N$14431 N$14528 N$14530 "Waveguide Crossing" sch_x=-112 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3769 N$14433 N$14435 N$14532 N$14534 "Waveguide Crossing" sch_x=-112 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3770 N$14437 N$14439 N$14536 N$14538 "Waveguide Crossing" sch_x=-112 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3771 N$14441 N$14443 N$14540 N$14542 "Waveguide Crossing" sch_x=-112 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3772 N$14445 N$14447 N$14544 N$14546 "Waveguide Crossing" sch_x=-112 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3773 N$14449 N$14451 N$14548 N$14550 "Waveguide Crossing" sch_x=-112 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3774 N$14453 N$14455 N$14552 N$14554 "Waveguide Crossing" sch_x=-112 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3775 N$14457 N$14459 N$14556 N$14558 "Waveguide Crossing" sch_x=-112 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3776 N$14461 N$14463 N$14560 N$14562 "Waveguide Crossing" sch_x=-112 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3777 N$14465 N$14467 N$14564 N$14566 "Waveguide Crossing" sch_x=-112 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3778 N$14469 N$14471 N$14568 N$14570 "Waveguide Crossing" sch_x=-112 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3779 N$14473 N$14475 N$14572 N$14574 "Waveguide Crossing" sch_x=-112 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3780 N$14477 N$14479 N$14576 N$15791 "Waveguide Crossing" sch_x=-112 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3781 N$14481 N$14483 N$15695 N$14578 "Waveguide Crossing" sch_x=-110 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3782 N$14485 N$14487 N$14580 N$14582 "Waveguide Crossing" sch_x=-110 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3783 N$14489 N$14491 N$14584 N$14586 "Waveguide Crossing" sch_x=-110 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3784 N$14493 N$14495 N$14588 N$14590 "Waveguide Crossing" sch_x=-110 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3785 N$14497 N$14499 N$14592 N$14594 "Waveguide Crossing" sch_x=-110 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3786 N$14501 N$14503 N$14596 N$14598 "Waveguide Crossing" sch_x=-110 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3787 N$14505 N$14507 N$14600 N$14602 "Waveguide Crossing" sch_x=-110 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3788 N$14509 N$14511 N$14604 N$14606 "Waveguide Crossing" sch_x=-110 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3789 N$14513 N$14515 N$14608 N$14610 "Waveguide Crossing" sch_x=-110 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3790 N$14517 N$14519 N$14612 N$14614 "Waveguide Crossing" sch_x=-110 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3791 N$14521 N$14523 N$14616 N$14618 "Waveguide Crossing" sch_x=-110 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3792 N$14525 N$14527 N$14620 N$14622 "Waveguide Crossing" sch_x=-110 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3793 N$14529 N$14531 N$14624 N$14626 "Waveguide Crossing" sch_x=-110 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3794 N$14533 N$14535 N$14628 N$14630 "Waveguide Crossing" sch_x=-110 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3795 N$14537 N$14539 N$14632 N$14634 "Waveguide Crossing" sch_x=-110 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3796 N$14541 N$14543 N$14636 N$14638 "Waveguide Crossing" sch_x=-110 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3797 N$14545 N$14547 N$14640 N$14642 "Waveguide Crossing" sch_x=-110 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3798 N$14549 N$14551 N$14644 N$14646 "Waveguide Crossing" sch_x=-110 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3799 N$14553 N$14555 N$14648 N$14650 "Waveguide Crossing" sch_x=-110 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3800 N$14557 N$14559 N$14652 N$14654 "Waveguide Crossing" sch_x=-110 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3801 N$14561 N$14563 N$14656 N$14658 "Waveguide Crossing" sch_x=-110 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3802 N$14565 N$14567 N$14660 N$14662 "Waveguide Crossing" sch_x=-110 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3803 N$14569 N$14571 N$14664 N$14666 "Waveguide Crossing" sch_x=-110 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3804 N$14573 N$14575 N$14668 N$15789 "Waveguide Crossing" sch_x=-110 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3805 N$14577 N$14579 N$15697 N$14670 "Waveguide Crossing" sch_x=-108 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3806 N$14581 N$14583 N$14672 N$14674 "Waveguide Crossing" sch_x=-108 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3807 N$14585 N$14587 N$14676 N$14678 "Waveguide Crossing" sch_x=-108 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3808 N$14589 N$14591 N$14680 N$14682 "Waveguide Crossing" sch_x=-108 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3809 N$14593 N$14595 N$14684 N$14686 "Waveguide Crossing" sch_x=-108 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3810 N$14597 N$14599 N$14688 N$14690 "Waveguide Crossing" sch_x=-108 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3811 N$14601 N$14603 N$14692 N$14694 "Waveguide Crossing" sch_x=-108 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3812 N$14605 N$14607 N$14696 N$14698 "Waveguide Crossing" sch_x=-108 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3813 N$14609 N$14611 N$14700 N$14702 "Waveguide Crossing" sch_x=-108 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3814 N$14613 N$14615 N$14704 N$14706 "Waveguide Crossing" sch_x=-108 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3815 N$14617 N$14619 N$14708 N$14710 "Waveguide Crossing" sch_x=-108 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3816 N$14621 N$14623 N$14712 N$14714 "Waveguide Crossing" sch_x=-108 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3817 N$14625 N$14627 N$14716 N$14718 "Waveguide Crossing" sch_x=-108 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3818 N$14629 N$14631 N$14720 N$14722 "Waveguide Crossing" sch_x=-108 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3819 N$14633 N$14635 N$14724 N$14726 "Waveguide Crossing" sch_x=-108 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3820 N$14637 N$14639 N$14728 N$14730 "Waveguide Crossing" sch_x=-108 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3821 N$14641 N$14643 N$14732 N$14734 "Waveguide Crossing" sch_x=-108 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3822 N$14645 N$14647 N$14736 N$14738 "Waveguide Crossing" sch_x=-108 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3823 N$14649 N$14651 N$14740 N$14742 "Waveguide Crossing" sch_x=-108 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3824 N$14653 N$14655 N$14744 N$14746 "Waveguide Crossing" sch_x=-108 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3825 N$14657 N$14659 N$14748 N$14750 "Waveguide Crossing" sch_x=-108 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3826 N$14661 N$14663 N$14752 N$14754 "Waveguide Crossing" sch_x=-108 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3827 N$14665 N$14667 N$14756 N$15787 "Waveguide Crossing" sch_x=-108 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3828 N$14669 N$14671 N$15699 N$14758 "Waveguide Crossing" sch_x=-106 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3829 N$14673 N$14675 N$14760 N$14762 "Waveguide Crossing" sch_x=-106 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3830 N$14677 N$14679 N$14764 N$14766 "Waveguide Crossing" sch_x=-106 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3831 N$14681 N$14683 N$14768 N$14770 "Waveguide Crossing" sch_x=-106 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3832 N$14685 N$14687 N$14772 N$14774 "Waveguide Crossing" sch_x=-106 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3833 N$14689 N$14691 N$14776 N$14778 "Waveguide Crossing" sch_x=-106 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3834 N$14693 N$14695 N$14780 N$14782 "Waveguide Crossing" sch_x=-106 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3835 N$14697 N$14699 N$14784 N$14786 "Waveguide Crossing" sch_x=-106 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3836 N$14701 N$14703 N$14788 N$14790 "Waveguide Crossing" sch_x=-106 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3837 N$14705 N$14707 N$14792 N$14794 "Waveguide Crossing" sch_x=-106 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3838 N$14709 N$14711 N$14796 N$14798 "Waveguide Crossing" sch_x=-106 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3839 N$14713 N$14715 N$14800 N$14802 "Waveguide Crossing" sch_x=-106 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3840 N$14717 N$14719 N$14804 N$14806 "Waveguide Crossing" sch_x=-106 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3841 N$14721 N$14723 N$14808 N$14810 "Waveguide Crossing" sch_x=-106 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3842 N$14725 N$14727 N$14812 N$14814 "Waveguide Crossing" sch_x=-106 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3843 N$14729 N$14731 N$14816 N$14818 "Waveguide Crossing" sch_x=-106 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3844 N$14733 N$14735 N$14820 N$14822 "Waveguide Crossing" sch_x=-106 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3845 N$14737 N$14739 N$14824 N$14826 "Waveguide Crossing" sch_x=-106 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3846 N$14741 N$14743 N$14828 N$14830 "Waveguide Crossing" sch_x=-106 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3847 N$14745 N$14747 N$14832 N$14834 "Waveguide Crossing" sch_x=-106 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3848 N$14749 N$14751 N$14836 N$14838 "Waveguide Crossing" sch_x=-106 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3849 N$14753 N$14755 N$14840 N$15785 "Waveguide Crossing" sch_x=-106 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3850 N$14757 N$14759 N$15701 N$14842 "Waveguide Crossing" sch_x=-104 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3851 N$14761 N$14763 N$14844 N$14846 "Waveguide Crossing" sch_x=-104 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3852 N$14765 N$14767 N$14848 N$14850 "Waveguide Crossing" sch_x=-104 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3853 N$14769 N$14771 N$14852 N$14854 "Waveguide Crossing" sch_x=-104 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3854 N$14773 N$14775 N$14856 N$14858 "Waveguide Crossing" sch_x=-104 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3855 N$14777 N$14779 N$14860 N$14862 "Waveguide Crossing" sch_x=-104 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3856 N$14781 N$14783 N$14864 N$14866 "Waveguide Crossing" sch_x=-104 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3857 N$14785 N$14787 N$14868 N$14870 "Waveguide Crossing" sch_x=-104 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3858 N$14789 N$14791 N$14872 N$14874 "Waveguide Crossing" sch_x=-104 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3859 N$14793 N$14795 N$14876 N$14878 "Waveguide Crossing" sch_x=-104 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3860 N$14797 N$14799 N$14880 N$14882 "Waveguide Crossing" sch_x=-104 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3861 N$14801 N$14803 N$14884 N$14886 "Waveguide Crossing" sch_x=-104 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3862 N$14805 N$14807 N$14888 N$14890 "Waveguide Crossing" sch_x=-104 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3863 N$14809 N$14811 N$14892 N$14894 "Waveguide Crossing" sch_x=-104 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3864 N$14813 N$14815 N$14896 N$14898 "Waveguide Crossing" sch_x=-104 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3865 N$14817 N$14819 N$14900 N$14902 "Waveguide Crossing" sch_x=-104 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3866 N$14821 N$14823 N$14904 N$14906 "Waveguide Crossing" sch_x=-104 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3867 N$14825 N$14827 N$14908 N$14910 "Waveguide Crossing" sch_x=-104 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3868 N$14829 N$14831 N$14912 N$14914 "Waveguide Crossing" sch_x=-104 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3869 N$14833 N$14835 N$14916 N$14918 "Waveguide Crossing" sch_x=-104 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3870 N$14837 N$14839 N$14920 N$15783 "Waveguide Crossing" sch_x=-104 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3871 N$14841 N$14843 N$15703 N$14922 "Waveguide Crossing" sch_x=-102 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3872 N$14845 N$14847 N$14924 N$14926 "Waveguide Crossing" sch_x=-102 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3873 N$14849 N$14851 N$14928 N$14930 "Waveguide Crossing" sch_x=-102 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3874 N$14853 N$14855 N$14932 N$14934 "Waveguide Crossing" sch_x=-102 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3875 N$14857 N$14859 N$14936 N$14938 "Waveguide Crossing" sch_x=-102 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3876 N$14861 N$14863 N$14940 N$14942 "Waveguide Crossing" sch_x=-102 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3877 N$14865 N$14867 N$14944 N$14946 "Waveguide Crossing" sch_x=-102 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3878 N$14869 N$14871 N$14948 N$14950 "Waveguide Crossing" sch_x=-102 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3879 N$14873 N$14875 N$14952 N$14954 "Waveguide Crossing" sch_x=-102 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3880 N$14877 N$14879 N$14956 N$14958 "Waveguide Crossing" sch_x=-102 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3881 N$14881 N$14883 N$14960 N$14962 "Waveguide Crossing" sch_x=-102 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3882 N$14885 N$14887 N$14964 N$14966 "Waveguide Crossing" sch_x=-102 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3883 N$14889 N$14891 N$14968 N$14970 "Waveguide Crossing" sch_x=-102 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3884 N$14893 N$14895 N$14972 N$14974 "Waveguide Crossing" sch_x=-102 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3885 N$14897 N$14899 N$14976 N$14978 "Waveguide Crossing" sch_x=-102 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3886 N$14901 N$14903 N$14980 N$14982 "Waveguide Crossing" sch_x=-102 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3887 N$14905 N$14907 N$14984 N$14986 "Waveguide Crossing" sch_x=-102 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3888 N$14909 N$14911 N$14988 N$14990 "Waveguide Crossing" sch_x=-102 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3889 N$14913 N$14915 N$14992 N$14994 "Waveguide Crossing" sch_x=-102 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3890 N$14917 N$14919 N$14996 N$15781 "Waveguide Crossing" sch_x=-102 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3891 N$14921 N$14923 N$15705 N$14998 "Waveguide Crossing" sch_x=-100 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3892 N$14925 N$14927 N$15000 N$15002 "Waveguide Crossing" sch_x=-100 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3893 N$14929 N$14931 N$15004 N$15006 "Waveguide Crossing" sch_x=-100 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3894 N$14933 N$14935 N$15008 N$15010 "Waveguide Crossing" sch_x=-100 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3895 N$14937 N$14939 N$15012 N$15014 "Waveguide Crossing" sch_x=-100 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3896 N$14941 N$14943 N$15016 N$15018 "Waveguide Crossing" sch_x=-100 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3897 N$14945 N$14947 N$15020 N$15022 "Waveguide Crossing" sch_x=-100 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3898 N$14949 N$14951 N$15024 N$15026 "Waveguide Crossing" sch_x=-100 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3899 N$14953 N$14955 N$15028 N$15030 "Waveguide Crossing" sch_x=-100 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3900 N$14957 N$14959 N$15032 N$15034 "Waveguide Crossing" sch_x=-100 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3901 N$14961 N$14963 N$15036 N$15038 "Waveguide Crossing" sch_x=-100 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3902 N$14965 N$14967 N$15040 N$15042 "Waveguide Crossing" sch_x=-100 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3903 N$14969 N$14971 N$15044 N$15046 "Waveguide Crossing" sch_x=-100 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3904 N$14973 N$14975 N$15048 N$15050 "Waveguide Crossing" sch_x=-100 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3905 N$14977 N$14979 N$15052 N$15054 "Waveguide Crossing" sch_x=-100 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3906 N$14981 N$14983 N$15056 N$15058 "Waveguide Crossing" sch_x=-100 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3907 N$14985 N$14987 N$15060 N$15062 "Waveguide Crossing" sch_x=-100 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3908 N$14989 N$14991 N$15064 N$15066 "Waveguide Crossing" sch_x=-100 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3909 N$14993 N$14995 N$15068 N$15779 "Waveguide Crossing" sch_x=-100 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3910 N$14997 N$14999 N$15707 N$15070 "Waveguide Crossing" sch_x=-98 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3911 N$15001 N$15003 N$15072 N$15074 "Waveguide Crossing" sch_x=-98 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3912 N$15005 N$15007 N$15076 N$15078 "Waveguide Crossing" sch_x=-98 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3913 N$15009 N$15011 N$15080 N$15082 "Waveguide Crossing" sch_x=-98 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3914 N$15013 N$15015 N$15084 N$15086 "Waveguide Crossing" sch_x=-98 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3915 N$15017 N$15019 N$15088 N$15090 "Waveguide Crossing" sch_x=-98 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3916 N$15021 N$15023 N$15092 N$15094 "Waveguide Crossing" sch_x=-98 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3917 N$15025 N$15027 N$15096 N$15098 "Waveguide Crossing" sch_x=-98 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3918 N$15029 N$15031 N$15100 N$15102 "Waveguide Crossing" sch_x=-98 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3919 N$15033 N$15035 N$15104 N$15106 "Waveguide Crossing" sch_x=-98 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3920 N$15037 N$15039 N$15108 N$15110 "Waveguide Crossing" sch_x=-98 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3921 N$15041 N$15043 N$15112 N$15114 "Waveguide Crossing" sch_x=-98 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3922 N$15045 N$15047 N$15116 N$15118 "Waveguide Crossing" sch_x=-98 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3923 N$15049 N$15051 N$15120 N$15122 "Waveguide Crossing" sch_x=-98 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3924 N$15053 N$15055 N$15124 N$15126 "Waveguide Crossing" sch_x=-98 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3925 N$15057 N$15059 N$15128 N$15130 "Waveguide Crossing" sch_x=-98 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3926 N$15061 N$15063 N$15132 N$15134 "Waveguide Crossing" sch_x=-98 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3927 N$15065 N$15067 N$15136 N$15777 "Waveguide Crossing" sch_x=-98 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3928 N$15069 N$15071 N$15709 N$15138 "Waveguide Crossing" sch_x=-96 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3929 N$15073 N$15075 N$15140 N$15142 "Waveguide Crossing" sch_x=-96 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3930 N$15077 N$15079 N$15144 N$15146 "Waveguide Crossing" sch_x=-96 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3931 N$15081 N$15083 N$15148 N$15150 "Waveguide Crossing" sch_x=-96 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3932 N$15085 N$15087 N$15152 N$15154 "Waveguide Crossing" sch_x=-96 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3933 N$15089 N$15091 N$15156 N$15158 "Waveguide Crossing" sch_x=-96 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3934 N$15093 N$15095 N$15160 N$15162 "Waveguide Crossing" sch_x=-96 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3935 N$15097 N$15099 N$15164 N$15166 "Waveguide Crossing" sch_x=-96 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3936 N$15101 N$15103 N$15168 N$15170 "Waveguide Crossing" sch_x=-96 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3937 N$15105 N$15107 N$15172 N$15174 "Waveguide Crossing" sch_x=-96 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3938 N$15109 N$15111 N$15176 N$15178 "Waveguide Crossing" sch_x=-96 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3939 N$15113 N$15115 N$15180 N$15182 "Waveguide Crossing" sch_x=-96 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3940 N$15117 N$15119 N$15184 N$15186 "Waveguide Crossing" sch_x=-96 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3941 N$15121 N$15123 N$15188 N$15190 "Waveguide Crossing" sch_x=-96 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3942 N$15125 N$15127 N$15192 N$15194 "Waveguide Crossing" sch_x=-96 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3943 N$15129 N$15131 N$15196 N$15198 "Waveguide Crossing" sch_x=-96 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3944 N$15133 N$15135 N$15200 N$15775 "Waveguide Crossing" sch_x=-96 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3945 N$15137 N$15139 N$15711 N$15202 "Waveguide Crossing" sch_x=-94 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3946 N$15141 N$15143 N$15204 N$15206 "Waveguide Crossing" sch_x=-94 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3947 N$15145 N$15147 N$15208 N$15210 "Waveguide Crossing" sch_x=-94 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3948 N$15149 N$15151 N$15212 N$15214 "Waveguide Crossing" sch_x=-94 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3949 N$15153 N$15155 N$15216 N$15218 "Waveguide Crossing" sch_x=-94 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3950 N$15157 N$15159 N$15220 N$15222 "Waveguide Crossing" sch_x=-94 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3951 N$15161 N$15163 N$15224 N$15226 "Waveguide Crossing" sch_x=-94 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3952 N$15165 N$15167 N$15228 N$15230 "Waveguide Crossing" sch_x=-94 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3953 N$15169 N$15171 N$15232 N$15234 "Waveguide Crossing" sch_x=-94 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3954 N$15173 N$15175 N$15236 N$15238 "Waveguide Crossing" sch_x=-94 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3955 N$15177 N$15179 N$15240 N$15242 "Waveguide Crossing" sch_x=-94 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3956 N$15181 N$15183 N$15244 N$15246 "Waveguide Crossing" sch_x=-94 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3957 N$15185 N$15187 N$15248 N$15250 "Waveguide Crossing" sch_x=-94 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3958 N$15189 N$15191 N$15252 N$15254 "Waveguide Crossing" sch_x=-94 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3959 N$15193 N$15195 N$15256 N$15258 "Waveguide Crossing" sch_x=-94 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3960 N$15197 N$15199 N$15260 N$15773 "Waveguide Crossing" sch_x=-94 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3961 N$15201 N$15203 N$15713 N$15262 "Waveguide Crossing" sch_x=-92 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3962 N$15205 N$15207 N$15264 N$15266 "Waveguide Crossing" sch_x=-92 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3963 N$15209 N$15211 N$15268 N$15270 "Waveguide Crossing" sch_x=-92 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3964 N$15213 N$15215 N$15272 N$15274 "Waveguide Crossing" sch_x=-92 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3965 N$15217 N$15219 N$15276 N$15278 "Waveguide Crossing" sch_x=-92 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3966 N$15221 N$15223 N$15280 N$15282 "Waveguide Crossing" sch_x=-92 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3967 N$15225 N$15227 N$15284 N$15286 "Waveguide Crossing" sch_x=-92 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3968 N$15229 N$15231 N$15288 N$15290 "Waveguide Crossing" sch_x=-92 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3969 N$15233 N$15235 N$15292 N$15294 "Waveguide Crossing" sch_x=-92 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3970 N$15237 N$15239 N$15296 N$15298 "Waveguide Crossing" sch_x=-92 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3971 N$15241 N$15243 N$15300 N$15302 "Waveguide Crossing" sch_x=-92 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3972 N$15245 N$15247 N$15304 N$15306 "Waveguide Crossing" sch_x=-92 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3973 N$15249 N$15251 N$15308 N$15310 "Waveguide Crossing" sch_x=-92 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3974 N$15253 N$15255 N$15312 N$15314 "Waveguide Crossing" sch_x=-92 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3975 N$15257 N$15259 N$15316 N$15771 "Waveguide Crossing" sch_x=-92 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3976 N$15261 N$15263 N$15715 N$15318 "Waveguide Crossing" sch_x=-90 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3977 N$15265 N$15267 N$15320 N$15322 "Waveguide Crossing" sch_x=-90 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3978 N$15269 N$15271 N$15324 N$15326 "Waveguide Crossing" sch_x=-90 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3979 N$15273 N$15275 N$15328 N$15330 "Waveguide Crossing" sch_x=-90 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3980 N$15277 N$15279 N$15332 N$15334 "Waveguide Crossing" sch_x=-90 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3981 N$15281 N$15283 N$15336 N$15338 "Waveguide Crossing" sch_x=-90 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3982 N$15285 N$15287 N$15340 N$15342 "Waveguide Crossing" sch_x=-90 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3983 N$15289 N$15291 N$15344 N$15346 "Waveguide Crossing" sch_x=-90 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3984 N$15293 N$15295 N$15348 N$15350 "Waveguide Crossing" sch_x=-90 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3985 N$15297 N$15299 N$15352 N$15354 "Waveguide Crossing" sch_x=-90 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3986 N$15301 N$15303 N$15356 N$15358 "Waveguide Crossing" sch_x=-90 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3987 N$15305 N$15307 N$15360 N$15362 "Waveguide Crossing" sch_x=-90 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3988 N$15309 N$15311 N$15364 N$15366 "Waveguide Crossing" sch_x=-90 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3989 N$15313 N$15315 N$15368 N$15769 "Waveguide Crossing" sch_x=-90 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3990 N$15317 N$15319 N$15717 N$15370 "Waveguide Crossing" sch_x=-88 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3991 N$15321 N$15323 N$15372 N$15374 "Waveguide Crossing" sch_x=-88 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3992 N$15325 N$15327 N$15376 N$15378 "Waveguide Crossing" sch_x=-88 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3993 N$15329 N$15331 N$15380 N$15382 "Waveguide Crossing" sch_x=-88 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3994 N$15333 N$15335 N$15384 N$15386 "Waveguide Crossing" sch_x=-88 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3995 N$15337 N$15339 N$15388 N$15390 "Waveguide Crossing" sch_x=-88 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3996 N$15341 N$15343 N$15392 N$15394 "Waveguide Crossing" sch_x=-88 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3997 N$15345 N$15347 N$15396 N$15398 "Waveguide Crossing" sch_x=-88 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3998 N$15349 N$15351 N$15400 N$15402 "Waveguide Crossing" sch_x=-88 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3999 N$15353 N$15355 N$15404 N$15406 "Waveguide Crossing" sch_x=-88 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4000 N$15357 N$15359 N$15408 N$15410 "Waveguide Crossing" sch_x=-88 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4001 N$15361 N$15363 N$15412 N$15414 "Waveguide Crossing" sch_x=-88 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4002 N$15365 N$15367 N$15416 N$15767 "Waveguide Crossing" sch_x=-88 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4003 N$15369 N$15371 N$15719 N$15418 "Waveguide Crossing" sch_x=-86 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4004 N$15373 N$15375 N$15420 N$15422 "Waveguide Crossing" sch_x=-86 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4005 N$15377 N$15379 N$15424 N$15426 "Waveguide Crossing" sch_x=-86 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4006 N$15381 N$15383 N$15428 N$15430 "Waveguide Crossing" sch_x=-86 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4007 N$15385 N$15387 N$15432 N$15434 "Waveguide Crossing" sch_x=-86 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4008 N$15389 N$15391 N$15436 N$15438 "Waveguide Crossing" sch_x=-86 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4009 N$15393 N$15395 N$15440 N$15442 "Waveguide Crossing" sch_x=-86 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4010 N$15397 N$15399 N$15444 N$15446 "Waveguide Crossing" sch_x=-86 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4011 N$15401 N$15403 N$15448 N$15450 "Waveguide Crossing" sch_x=-86 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4012 N$15405 N$15407 N$15452 N$15454 "Waveguide Crossing" sch_x=-86 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4013 N$15409 N$15411 N$15456 N$15458 "Waveguide Crossing" sch_x=-86 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4014 N$15413 N$15415 N$15460 N$15765 "Waveguide Crossing" sch_x=-86 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4015 N$15417 N$15419 N$15721 N$15462 "Waveguide Crossing" sch_x=-84 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4016 N$15421 N$15423 N$15464 N$15466 "Waveguide Crossing" sch_x=-84 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4017 N$15425 N$15427 N$15468 N$15470 "Waveguide Crossing" sch_x=-84 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4018 N$15429 N$15431 N$15472 N$15474 "Waveguide Crossing" sch_x=-84 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4019 N$15433 N$15435 N$15476 N$15478 "Waveguide Crossing" sch_x=-84 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4020 N$15437 N$15439 N$15480 N$15482 "Waveguide Crossing" sch_x=-84 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4021 N$15441 N$15443 N$15484 N$15486 "Waveguide Crossing" sch_x=-84 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4022 N$15445 N$15447 N$15488 N$15490 "Waveguide Crossing" sch_x=-84 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4023 N$15449 N$15451 N$15492 N$15494 "Waveguide Crossing" sch_x=-84 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4024 N$15453 N$15455 N$15496 N$15498 "Waveguide Crossing" sch_x=-84 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4025 N$15457 N$15459 N$15500 N$15763 "Waveguide Crossing" sch_x=-84 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4026 N$15461 N$15463 N$15723 N$15502 "Waveguide Crossing" sch_x=-82 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4027 N$15465 N$15467 N$15504 N$15506 "Waveguide Crossing" sch_x=-82 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4028 N$15469 N$15471 N$15508 N$15510 "Waveguide Crossing" sch_x=-82 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4029 N$15473 N$15475 N$15512 N$15514 "Waveguide Crossing" sch_x=-82 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4030 N$15477 N$15479 N$15516 N$15518 "Waveguide Crossing" sch_x=-82 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4031 N$15481 N$15483 N$15520 N$15522 "Waveguide Crossing" sch_x=-82 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4032 N$15485 N$15487 N$15524 N$15526 "Waveguide Crossing" sch_x=-82 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4033 N$15489 N$15491 N$15528 N$15530 "Waveguide Crossing" sch_x=-82 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4034 N$15493 N$15495 N$15532 N$15534 "Waveguide Crossing" sch_x=-82 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4035 N$15497 N$15499 N$15536 N$15761 "Waveguide Crossing" sch_x=-82 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4036 N$15501 N$15503 N$15725 N$15538 "Waveguide Crossing" sch_x=-80 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4037 N$15505 N$15507 N$15540 N$15542 "Waveguide Crossing" sch_x=-80 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4038 N$15509 N$15511 N$15544 N$15546 "Waveguide Crossing" sch_x=-80 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4039 N$15513 N$15515 N$15548 N$15550 "Waveguide Crossing" sch_x=-80 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4040 N$15517 N$15519 N$15552 N$15554 "Waveguide Crossing" sch_x=-80 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4041 N$15521 N$15523 N$15556 N$15558 "Waveguide Crossing" sch_x=-80 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4042 N$15525 N$15527 N$15560 N$15562 "Waveguide Crossing" sch_x=-80 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4043 N$15529 N$15531 N$15564 N$15566 "Waveguide Crossing" sch_x=-80 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4044 N$15533 N$15535 N$15568 N$15759 "Waveguide Crossing" sch_x=-80 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4045 N$15537 N$15539 N$15727 N$15570 "Waveguide Crossing" sch_x=-78 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4046 N$15541 N$15543 N$15572 N$15574 "Waveguide Crossing" sch_x=-78 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4047 N$15545 N$15547 N$15576 N$15578 "Waveguide Crossing" sch_x=-78 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4048 N$15549 N$15551 N$15580 N$15582 "Waveguide Crossing" sch_x=-78 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4049 N$15553 N$15555 N$15584 N$15586 "Waveguide Crossing" sch_x=-78 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4050 N$15557 N$15559 N$15588 N$15590 "Waveguide Crossing" sch_x=-78 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4051 N$15561 N$15563 N$15592 N$15594 "Waveguide Crossing" sch_x=-78 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4052 N$15565 N$15567 N$15596 N$15757 "Waveguide Crossing" sch_x=-78 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4053 N$15569 N$15571 N$15729 N$15598 "Waveguide Crossing" sch_x=-76 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4054 N$15573 N$15575 N$15600 N$15602 "Waveguide Crossing" sch_x=-76 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4055 N$15577 N$15579 N$15604 N$15606 "Waveguide Crossing" sch_x=-76 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4056 N$15581 N$15583 N$15608 N$15610 "Waveguide Crossing" sch_x=-76 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4057 N$15585 N$15587 N$15612 N$15614 "Waveguide Crossing" sch_x=-76 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4058 N$15589 N$15591 N$15616 N$15618 "Waveguide Crossing" sch_x=-76 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4059 N$15593 N$15595 N$15620 N$15755 "Waveguide Crossing" sch_x=-76 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4060 N$15597 N$15599 N$15731 N$15622 "Waveguide Crossing" sch_x=-74 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4061 N$15601 N$15603 N$15624 N$15626 "Waveguide Crossing" sch_x=-74 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4062 N$15605 N$15607 N$15628 N$15630 "Waveguide Crossing" sch_x=-74 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4063 N$15609 N$15611 N$15632 N$15634 "Waveguide Crossing" sch_x=-74 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4064 N$15613 N$15615 N$15636 N$15638 "Waveguide Crossing" sch_x=-74 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4065 N$15617 N$15619 N$15640 N$15753 "Waveguide Crossing" sch_x=-74 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4066 N$15621 N$15623 N$15733 N$15642 "Waveguide Crossing" sch_x=-72 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4067 N$15625 N$15627 N$15644 N$15646 "Waveguide Crossing" sch_x=-72 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4068 N$15629 N$15631 N$15648 N$15650 "Waveguide Crossing" sch_x=-72 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4069 N$15633 N$15635 N$15652 N$15654 "Waveguide Crossing" sch_x=-72 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4070 N$15637 N$15639 N$15656 N$15751 "Waveguide Crossing" sch_x=-72 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4071 N$15641 N$15643 N$15735 N$15658 "Waveguide Crossing" sch_x=-70 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4072 N$15645 N$15647 N$15660 N$15662 "Waveguide Crossing" sch_x=-70 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4073 N$15649 N$15651 N$15664 N$15666 "Waveguide Crossing" sch_x=-70 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4074 N$15653 N$15655 N$15668 N$15749 "Waveguide Crossing" sch_x=-70 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4075 N$15657 N$15659 N$15737 N$15670 "Waveguide Crossing" sch_x=-68 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4076 N$15661 N$15663 N$15672 N$15674 "Waveguide Crossing" sch_x=-68 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4077 N$15665 N$15667 N$15676 N$15747 "Waveguide Crossing" sch_x=-68 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4078 N$15669 N$15671 N$15739 N$15678 "Waveguide Crossing" sch_x=-66 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4079 N$15673 N$15675 N$15680 N$15745 "Waveguide Crossing" sch_x=-66 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4080 N$15677 N$15679 N$15741 N$15743 "Waveguide Crossing" sch_x=-64 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3281 N$15744 N$15746 N$13149 N$12610 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3282 N$15748 N$15750 N$12612 N$12614 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3283 N$15752 N$15754 N$12616 N$12618 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3284 N$15756 N$15758 N$12620 N$12622 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3285 N$15760 N$15762 N$12624 N$12626 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3286 N$15764 N$15766 N$12628 N$12630 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3287 N$15768 N$15770 N$12632 N$12634 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3288 N$15772 N$15774 N$12636 N$12638 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3289 N$15776 N$15778 N$12640 N$12642 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3290 N$15780 N$15782 N$12644 N$12646 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3291 N$15784 N$15786 N$12648 N$12650 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3292 N$15788 N$15790 N$12652 N$12654 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3293 N$15792 N$15794 N$12656 N$12658 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3294 N$15796 N$15798 N$12660 N$12662 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3295 N$15800 N$15802 N$12664 N$12666 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3296 N$15804 N$15808 N$12668 N$13151 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3297 N$12609 N$12611 N$13089 N$12670 "Waveguide Crossing" sch_x=-60 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3298 N$12613 N$12615 N$12672 N$12674 "Waveguide Crossing" sch_x=-60 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3299 N$12617 N$12619 N$12676 N$12678 "Waveguide Crossing" sch_x=-60 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3300 N$12621 N$12623 N$12680 N$12682 "Waveguide Crossing" sch_x=-60 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3301 N$12625 N$12627 N$12684 N$12686 "Waveguide Crossing" sch_x=-60 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3302 N$12629 N$12631 N$12688 N$12690 "Waveguide Crossing" sch_x=-60 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3303 N$12633 N$12635 N$12692 N$12694 "Waveguide Crossing" sch_x=-60 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3304 N$12637 N$12639 N$12696 N$12698 "Waveguide Crossing" sch_x=-60 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3305 N$12641 N$12643 N$12700 N$12702 "Waveguide Crossing" sch_x=-60 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3306 N$12645 N$12647 N$12704 N$12706 "Waveguide Crossing" sch_x=-60 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3307 N$12649 N$12651 N$12708 N$12710 "Waveguide Crossing" sch_x=-60 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3308 N$12653 N$12655 N$12712 N$12714 "Waveguide Crossing" sch_x=-60 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3309 N$12657 N$12659 N$12716 N$12718 "Waveguide Crossing" sch_x=-60 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3310 N$12661 N$12663 N$12720 N$12722 "Waveguide Crossing" sch_x=-60 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3311 N$12665 N$12667 N$12724 N$13147 "Waveguide Crossing" sch_x=-60 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3312 N$12669 N$12671 N$13091 N$12726 "Waveguide Crossing" sch_x=-58 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3313 N$12673 N$12675 N$12728 N$12730 "Waveguide Crossing" sch_x=-58 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3314 N$12677 N$12679 N$12732 N$12734 "Waveguide Crossing" sch_x=-58 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3315 N$12681 N$12683 N$12736 N$12738 "Waveguide Crossing" sch_x=-58 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3316 N$12685 N$12687 N$12740 N$12742 "Waveguide Crossing" sch_x=-58 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3317 N$12689 N$12691 N$12744 N$12746 "Waveguide Crossing" sch_x=-58 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3318 N$12693 N$12695 N$12748 N$12750 "Waveguide Crossing" sch_x=-58 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3319 N$12697 N$12699 N$12752 N$12754 "Waveguide Crossing" sch_x=-58 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3320 N$12701 N$12703 N$12756 N$12758 "Waveguide Crossing" sch_x=-58 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3321 N$12705 N$12707 N$12760 N$12762 "Waveguide Crossing" sch_x=-58 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3322 N$12709 N$12711 N$12764 N$12766 "Waveguide Crossing" sch_x=-58 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3323 N$12713 N$12715 N$12768 N$12770 "Waveguide Crossing" sch_x=-58 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3324 N$12717 N$12719 N$12772 N$12774 "Waveguide Crossing" sch_x=-58 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3325 N$12721 N$12723 N$12776 N$13145 "Waveguide Crossing" sch_x=-58 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3326 N$12725 N$12727 N$13093 N$12778 "Waveguide Crossing" sch_x=-56 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3327 N$12729 N$12731 N$12780 N$12782 "Waveguide Crossing" sch_x=-56 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3328 N$12733 N$12735 N$12784 N$12786 "Waveguide Crossing" sch_x=-56 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3329 N$12737 N$12739 N$12788 N$12790 "Waveguide Crossing" sch_x=-56 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3330 N$12741 N$12743 N$12792 N$12794 "Waveguide Crossing" sch_x=-56 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3331 N$12745 N$12747 N$12796 N$12798 "Waveguide Crossing" sch_x=-56 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3332 N$12749 N$12751 N$12800 N$12802 "Waveguide Crossing" sch_x=-56 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3333 N$12753 N$12755 N$12804 N$12806 "Waveguide Crossing" sch_x=-56 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3334 N$12757 N$12759 N$12808 N$12810 "Waveguide Crossing" sch_x=-56 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3335 N$12761 N$12763 N$12812 N$12814 "Waveguide Crossing" sch_x=-56 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3336 N$12765 N$12767 N$12816 N$12818 "Waveguide Crossing" sch_x=-56 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3337 N$12769 N$12771 N$12820 N$12822 "Waveguide Crossing" sch_x=-56 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3338 N$12773 N$12775 N$12824 N$13143 "Waveguide Crossing" sch_x=-56 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3339 N$12777 N$12779 N$13095 N$12826 "Waveguide Crossing" sch_x=-54 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3340 N$12781 N$12783 N$12828 N$12830 "Waveguide Crossing" sch_x=-54 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3341 N$12785 N$12787 N$12832 N$12834 "Waveguide Crossing" sch_x=-54 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3342 N$12789 N$12791 N$12836 N$12838 "Waveguide Crossing" sch_x=-54 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3343 N$12793 N$12795 N$12840 N$12842 "Waveguide Crossing" sch_x=-54 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3344 N$12797 N$12799 N$12844 N$12846 "Waveguide Crossing" sch_x=-54 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3345 N$12801 N$12803 N$12848 N$12850 "Waveguide Crossing" sch_x=-54 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3346 N$12805 N$12807 N$12852 N$12854 "Waveguide Crossing" sch_x=-54 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3347 N$12809 N$12811 N$12856 N$12858 "Waveguide Crossing" sch_x=-54 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3348 N$12813 N$12815 N$12860 N$12862 "Waveguide Crossing" sch_x=-54 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3349 N$12817 N$12819 N$12864 N$12866 "Waveguide Crossing" sch_x=-54 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3350 N$12821 N$12823 N$12868 N$13141 "Waveguide Crossing" sch_x=-54 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3351 N$12825 N$12827 N$13097 N$12870 "Waveguide Crossing" sch_x=-52 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3352 N$12829 N$12831 N$12872 N$12874 "Waveguide Crossing" sch_x=-52 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3353 N$12833 N$12835 N$12876 N$12878 "Waveguide Crossing" sch_x=-52 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3354 N$12837 N$12839 N$12880 N$12882 "Waveguide Crossing" sch_x=-52 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3355 N$12841 N$12843 N$12884 N$12886 "Waveguide Crossing" sch_x=-52 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3356 N$12845 N$12847 N$12888 N$12890 "Waveguide Crossing" sch_x=-52 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3357 N$12849 N$12851 N$12892 N$12894 "Waveguide Crossing" sch_x=-52 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3358 N$12853 N$12855 N$12896 N$12898 "Waveguide Crossing" sch_x=-52 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3359 N$12857 N$12859 N$12900 N$12902 "Waveguide Crossing" sch_x=-52 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3360 N$12861 N$12863 N$12904 N$12906 "Waveguide Crossing" sch_x=-52 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3361 N$12865 N$12867 N$12908 N$13139 "Waveguide Crossing" sch_x=-52 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3362 N$12869 N$12871 N$13099 N$12910 "Waveguide Crossing" sch_x=-50 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3363 N$12873 N$12875 N$12912 N$12914 "Waveguide Crossing" sch_x=-50 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3364 N$12877 N$12879 N$12916 N$12918 "Waveguide Crossing" sch_x=-50 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3365 N$12881 N$12883 N$12920 N$12922 "Waveguide Crossing" sch_x=-50 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3366 N$12885 N$12887 N$12924 N$12926 "Waveguide Crossing" sch_x=-50 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3367 N$12889 N$12891 N$12928 N$12930 "Waveguide Crossing" sch_x=-50 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3368 N$12893 N$12895 N$12932 N$12934 "Waveguide Crossing" sch_x=-50 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3369 N$12897 N$12899 N$12936 N$12938 "Waveguide Crossing" sch_x=-50 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3370 N$12901 N$12903 N$12940 N$12942 "Waveguide Crossing" sch_x=-50 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3371 N$12905 N$12907 N$12944 N$13137 "Waveguide Crossing" sch_x=-50 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3372 N$12909 N$12911 N$13101 N$12946 "Waveguide Crossing" sch_x=-48 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3373 N$12913 N$12915 N$12948 N$12950 "Waveguide Crossing" sch_x=-48 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3374 N$12917 N$12919 N$12952 N$12954 "Waveguide Crossing" sch_x=-48 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3375 N$12921 N$12923 N$12956 N$12958 "Waveguide Crossing" sch_x=-48 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3376 N$12925 N$12927 N$12960 N$12962 "Waveguide Crossing" sch_x=-48 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3377 N$12929 N$12931 N$12964 N$12966 "Waveguide Crossing" sch_x=-48 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3378 N$12933 N$12935 N$12968 N$12970 "Waveguide Crossing" sch_x=-48 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3379 N$12937 N$12939 N$12972 N$12974 "Waveguide Crossing" sch_x=-48 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3380 N$12941 N$12943 N$12976 N$13135 "Waveguide Crossing" sch_x=-48 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3381 N$12945 N$12947 N$13103 N$12978 "Waveguide Crossing" sch_x=-46 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3382 N$12949 N$12951 N$12980 N$12982 "Waveguide Crossing" sch_x=-46 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3383 N$12953 N$12955 N$12984 N$12986 "Waveguide Crossing" sch_x=-46 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3384 N$12957 N$12959 N$12988 N$12990 "Waveguide Crossing" sch_x=-46 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3385 N$12961 N$12963 N$12992 N$12994 "Waveguide Crossing" sch_x=-46 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3386 N$12965 N$12967 N$12996 N$12998 "Waveguide Crossing" sch_x=-46 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3387 N$12969 N$12971 N$13000 N$13002 "Waveguide Crossing" sch_x=-46 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3388 N$12973 N$12975 N$13004 N$13133 "Waveguide Crossing" sch_x=-46 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3389 N$12977 N$12979 N$13105 N$13006 "Waveguide Crossing" sch_x=-44 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3390 N$12981 N$12983 N$13008 N$13010 "Waveguide Crossing" sch_x=-44 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3391 N$12985 N$12987 N$13012 N$13014 "Waveguide Crossing" sch_x=-44 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3392 N$12989 N$12991 N$13016 N$13018 "Waveguide Crossing" sch_x=-44 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3393 N$12993 N$12995 N$13020 N$13022 "Waveguide Crossing" sch_x=-44 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3394 N$12997 N$12999 N$13024 N$13026 "Waveguide Crossing" sch_x=-44 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3395 N$13001 N$13003 N$13028 N$13131 "Waveguide Crossing" sch_x=-44 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3396 N$13005 N$13007 N$13107 N$13030 "Waveguide Crossing" sch_x=-42 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3397 N$13009 N$13011 N$13032 N$13034 "Waveguide Crossing" sch_x=-42 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3398 N$13013 N$13015 N$13036 N$13038 "Waveguide Crossing" sch_x=-42 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3399 N$13017 N$13019 N$13040 N$13042 "Waveguide Crossing" sch_x=-42 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3400 N$13021 N$13023 N$13044 N$13046 "Waveguide Crossing" sch_x=-42 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3401 N$13025 N$13027 N$13048 N$13129 "Waveguide Crossing" sch_x=-42 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3402 N$13029 N$13031 N$13109 N$13050 "Waveguide Crossing" sch_x=-40 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3403 N$13033 N$13035 N$13052 N$13054 "Waveguide Crossing" sch_x=-40 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3404 N$13037 N$13039 N$13056 N$13058 "Waveguide Crossing" sch_x=-40 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3405 N$13041 N$13043 N$13060 N$13062 "Waveguide Crossing" sch_x=-40 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3406 N$13045 N$13047 N$13064 N$13127 "Waveguide Crossing" sch_x=-40 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3407 N$13049 N$13051 N$13111 N$13066 "Waveguide Crossing" sch_x=-38 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3408 N$13053 N$13055 N$13068 N$13070 "Waveguide Crossing" sch_x=-38 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3409 N$13057 N$13059 N$13072 N$13074 "Waveguide Crossing" sch_x=-38 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3410 N$13061 N$13063 N$13076 N$13125 "Waveguide Crossing" sch_x=-38 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3411 N$13065 N$13067 N$13113 N$13078 "Waveguide Crossing" sch_x=-36 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3412 N$13069 N$13071 N$13080 N$13082 "Waveguide Crossing" sch_x=-36 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3413 N$13073 N$13075 N$13084 N$13123 "Waveguide Crossing" sch_x=-36 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3414 N$13077 N$13079 N$13115 N$13086 "Waveguide Crossing" sch_x=-34 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3415 N$13081 N$13083 N$13088 N$13121 "Waveguide Crossing" sch_x=-34 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3416 N$13085 N$13087 N$13117 N$13119 "Waveguide Crossing" sch_x=-32 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3209 N$13120 N$13122 N$12461 N$12322 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3210 N$13124 N$13126 N$12324 N$12326 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3211 N$13128 N$13130 N$12328 N$12330 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3212 N$13132 N$13134 N$12332 N$12334 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3213 N$13136 N$13138 N$12336 N$12338 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3214 N$13140 N$13142 N$12340 N$12342 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3215 N$13144 N$13146 N$12344 N$12346 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3216 N$13148 N$13152 N$12348 N$12463 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3217 N$12321 N$12323 N$12433 N$12350 "Waveguide Crossing" sch_x=-28 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3218 N$12325 N$12327 N$12352 N$12354 "Waveguide Crossing" sch_x=-28 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3219 N$12329 N$12331 N$12356 N$12358 "Waveguide Crossing" sch_x=-28 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3220 N$12333 N$12335 N$12360 N$12362 "Waveguide Crossing" sch_x=-28 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3221 N$12337 N$12339 N$12364 N$12366 "Waveguide Crossing" sch_x=-28 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3222 N$12341 N$12343 N$12368 N$12370 "Waveguide Crossing" sch_x=-28 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3223 N$12345 N$12347 N$12372 N$12459 "Waveguide Crossing" sch_x=-28 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3224 N$12349 N$12351 N$12435 N$12374 "Waveguide Crossing" sch_x=-26 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3225 N$12353 N$12355 N$12376 N$12378 "Waveguide Crossing" sch_x=-26 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3226 N$12357 N$12359 N$12380 N$12382 "Waveguide Crossing" sch_x=-26 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3227 N$12361 N$12363 N$12384 N$12386 "Waveguide Crossing" sch_x=-26 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3228 N$12365 N$12367 N$12388 N$12390 "Waveguide Crossing" sch_x=-26 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3229 N$12369 N$12371 N$12392 N$12457 "Waveguide Crossing" sch_x=-26 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3230 N$12373 N$12375 N$12437 N$12394 "Waveguide Crossing" sch_x=-24 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3231 N$12377 N$12379 N$12396 N$12398 "Waveguide Crossing" sch_x=-24 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3232 N$12381 N$12383 N$12400 N$12402 "Waveguide Crossing" sch_x=-24 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3233 N$12385 N$12387 N$12404 N$12406 "Waveguide Crossing" sch_x=-24 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3234 N$12389 N$12391 N$12408 N$12455 "Waveguide Crossing" sch_x=-24 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3235 N$12393 N$12395 N$12439 N$12410 "Waveguide Crossing" sch_x=-22 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3236 N$12397 N$12399 N$12412 N$12414 "Waveguide Crossing" sch_x=-22 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3237 N$12401 N$12403 N$12416 N$12418 "Waveguide Crossing" sch_x=-22 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3238 N$12405 N$12407 N$12420 N$12453 "Waveguide Crossing" sch_x=-22 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3239 N$12409 N$12411 N$12441 N$12422 "Waveguide Crossing" sch_x=-20 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3240 N$12413 N$12415 N$12424 N$12426 "Waveguide Crossing" sch_x=-20 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3241 N$12417 N$12419 N$12428 N$12451 "Waveguide Crossing" sch_x=-20 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3242 N$12421 N$12423 N$12443 N$12430 "Waveguide Crossing" sch_x=-18 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3243 N$12425 N$12427 N$12432 N$12449 "Waveguide Crossing" sch_x=-18 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3244 N$12429 N$12431 N$12445 N$12447 "Waveguide Crossing" sch_x=-16 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3189 N$12448 N$12450 N$12277 N$12242 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3190 N$12452 N$12454 N$12244 N$12246 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3191 N$12456 N$12458 N$12248 N$12250 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3192 N$12460 N$12464 N$12252 N$12279 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3193 N$12241 N$12243 N$12265 N$12254 "Waveguide Crossing" sch_x=-12 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3194 N$12245 N$12247 N$12256 N$12258 "Waveguide Crossing" sch_x=-12 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3195 N$12249 N$12251 N$12260 N$12275 "Waveguide Crossing" sch_x=-12 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3196 N$12253 N$12255 N$12267 N$12262 "Waveguide Crossing" sch_x=-10 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3197 N$12257 N$12259 N$12264 N$12273 "Waveguide Crossing" sch_x=-10 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3198 N$12261 N$12263 N$12269 N$12271 "Waveguide Crossing" sch_x=-8 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3137 N$12462 N$12434 N$12101 N$12066 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3138 N$12436 N$12438 N$12068 N$12070 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3139 N$12440 N$12442 N$12072 N$12074 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3140 N$12444 N$12446 N$12076 N$12103 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3141 N$12065 N$12067 N$12089 N$12078 "Waveguide Crossing" sch_x=-12 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3142 N$12069 N$12071 N$12080 N$12082 "Waveguide Crossing" sch_x=-12 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3143 N$12073 N$12075 N$12084 N$12099 "Waveguide Crossing" sch_x=-12 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3144 N$12077 N$12079 N$12091 N$12086 "Waveguide Crossing" sch_x=-10 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3145 N$12081 N$12083 N$12088 N$12097 "Waveguide Crossing" sch_x=-10 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3146 N$12085 N$12087 N$12093 N$12095 "Waveguide Crossing" sch_x=-8 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3033 N$13150 N$13090 N$11821 N$11682 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3034 N$13092 N$13094 N$11684 N$11686 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3035 N$13096 N$13098 N$11688 N$11690 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3036 N$13100 N$13102 N$11692 N$11694 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3037 N$13104 N$13106 N$11696 N$11698 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3038 N$13108 N$13110 N$11700 N$11702 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3039 N$13112 N$13114 N$11704 N$11706 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3040 N$13116 N$13118 N$11708 N$11823 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3041 N$11681 N$11683 N$11793 N$11710 "Waveguide Crossing" sch_x=-28 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3042 N$11685 N$11687 N$11712 N$11714 "Waveguide Crossing" sch_x=-28 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3043 N$11689 N$11691 N$11716 N$11718 "Waveguide Crossing" sch_x=-28 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3044 N$11693 N$11695 N$11720 N$11722 "Waveguide Crossing" sch_x=-28 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3045 N$11697 N$11699 N$11724 N$11726 "Waveguide Crossing" sch_x=-28 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3046 N$11701 N$11703 N$11728 N$11730 "Waveguide Crossing" sch_x=-28 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3047 N$11705 N$11707 N$11732 N$11819 "Waveguide Crossing" sch_x=-28 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3048 N$11709 N$11711 N$11795 N$11734 "Waveguide Crossing" sch_x=-26 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3049 N$11713 N$11715 N$11736 N$11738 "Waveguide Crossing" sch_x=-26 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3050 N$11717 N$11719 N$11740 N$11742 "Waveguide Crossing" sch_x=-26 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3051 N$11721 N$11723 N$11744 N$11746 "Waveguide Crossing" sch_x=-26 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3052 N$11725 N$11727 N$11748 N$11750 "Waveguide Crossing" sch_x=-26 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3053 N$11729 N$11731 N$11752 N$11817 "Waveguide Crossing" sch_x=-26 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3054 N$11733 N$11735 N$11797 N$11754 "Waveguide Crossing" sch_x=-24 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3055 N$11737 N$11739 N$11756 N$11758 "Waveguide Crossing" sch_x=-24 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3056 N$11741 N$11743 N$11760 N$11762 "Waveguide Crossing" sch_x=-24 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3057 N$11745 N$11747 N$11764 N$11766 "Waveguide Crossing" sch_x=-24 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3058 N$11749 N$11751 N$11768 N$11815 "Waveguide Crossing" sch_x=-24 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3059 N$11753 N$11755 N$11799 N$11770 "Waveguide Crossing" sch_x=-22 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3060 N$11757 N$11759 N$11772 N$11774 "Waveguide Crossing" sch_x=-22 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3061 N$11761 N$11763 N$11776 N$11778 "Waveguide Crossing" sch_x=-22 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3062 N$11765 N$11767 N$11780 N$11813 "Waveguide Crossing" sch_x=-22 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3063 N$11769 N$11771 N$11801 N$11782 "Waveguide Crossing" sch_x=-20 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3064 N$11773 N$11775 N$11784 N$11786 "Waveguide Crossing" sch_x=-20 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3065 N$11777 N$11779 N$11788 N$11811 "Waveguide Crossing" sch_x=-20 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3066 N$11781 N$11783 N$11803 N$11790 "Waveguide Crossing" sch_x=-18 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3067 N$11785 N$11787 N$11792 N$11809 "Waveguide Crossing" sch_x=-18 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3068 N$11789 N$11791 N$11805 N$11807 "Waveguide Crossing" sch_x=-16 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3013 N$11808 N$11810 N$11637 N$11602 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3014 N$11812 N$11814 N$11604 N$11606 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3015 N$11816 N$11818 N$11608 N$11610 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3016 N$11820 N$11824 N$11612 N$11639 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3017 N$11601 N$11603 N$11625 N$11614 "Waveguide Crossing" sch_x=-12 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3018 N$11605 N$11607 N$11616 N$11618 "Waveguide Crossing" sch_x=-12 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3019 N$11609 N$11611 N$11620 N$11635 "Waveguide Crossing" sch_x=-12 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3020 N$11613 N$11615 N$11627 N$11622 "Waveguide Crossing" sch_x=-10 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3021 N$11617 N$11619 N$11624 N$11633 "Waveguide Crossing" sch_x=-10 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3022 N$11621 N$11623 N$11629 N$11631 "Waveguide Crossing" sch_x=-8 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2961 N$11822 N$11794 N$11461 N$11426 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2962 N$11796 N$11798 N$11428 N$11430 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2963 N$11800 N$11802 N$11432 N$11434 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2964 N$11804 N$11806 N$11436 N$11463 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2965 N$11425 N$11427 N$11449 N$11438 "Waveguide Crossing" sch_x=-12 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2966 N$11429 N$11431 N$11440 N$11442 "Waveguide Crossing" sch_x=-12 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2967 N$11433 N$11435 N$11444 N$11459 "Waveguide Crossing" sch_x=-12 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2968 N$11437 N$11439 N$11451 N$11446 "Waveguide Crossing" sch_x=-10 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2969 N$11441 N$11443 N$11448 N$11457 "Waveguide Crossing" sch_x=-10 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2970 N$11445 N$11447 N$11453 N$11455 "Waveguide Crossing" sch_x=-8 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2657 N$15806 N$15682 N$10781 N$10242 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2658 N$15684 N$15686 N$10244 N$10246 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2659 N$15688 N$15690 N$10248 N$10250 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2660 N$15692 N$15694 N$10252 N$10254 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2661 N$15696 N$15698 N$10256 N$10258 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2662 N$15700 N$15702 N$10260 N$10262 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2663 N$15704 N$15706 N$10264 N$10266 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2664 N$15708 N$15710 N$10268 N$10270 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2665 N$15712 N$15714 N$10272 N$10274 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2666 N$15716 N$15718 N$10276 N$10278 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2667 N$15720 N$15722 N$10280 N$10282 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2668 N$15724 N$15726 N$10284 N$10286 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2669 N$15728 N$15730 N$10288 N$10290 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2670 N$15732 N$15734 N$10292 N$10294 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2671 N$15736 N$15738 N$10296 N$10298 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2672 N$15740 N$15742 N$10300 N$10783 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2673 N$10241 N$10243 N$10721 N$10302 "Waveguide Crossing" sch_x=-60 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2674 N$10245 N$10247 N$10304 N$10306 "Waveguide Crossing" sch_x=-60 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2675 N$10249 N$10251 N$10308 N$10310 "Waveguide Crossing" sch_x=-60 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2676 N$10253 N$10255 N$10312 N$10314 "Waveguide Crossing" sch_x=-60 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2677 N$10257 N$10259 N$10316 N$10318 "Waveguide Crossing" sch_x=-60 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2678 N$10261 N$10263 N$10320 N$10322 "Waveguide Crossing" sch_x=-60 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2679 N$10265 N$10267 N$10324 N$10326 "Waveguide Crossing" sch_x=-60 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2680 N$10269 N$10271 N$10328 N$10330 "Waveguide Crossing" sch_x=-60 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2681 N$10273 N$10275 N$10332 N$10334 "Waveguide Crossing" sch_x=-60 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2682 N$10277 N$10279 N$10336 N$10338 "Waveguide Crossing" sch_x=-60 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2683 N$10281 N$10283 N$10340 N$10342 "Waveguide Crossing" sch_x=-60 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2684 N$10285 N$10287 N$10344 N$10346 "Waveguide Crossing" sch_x=-60 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2685 N$10289 N$10291 N$10348 N$10350 "Waveguide Crossing" sch_x=-60 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2686 N$10293 N$10295 N$10352 N$10354 "Waveguide Crossing" sch_x=-60 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2687 N$10297 N$10299 N$10356 N$10779 "Waveguide Crossing" sch_x=-60 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2688 N$10301 N$10303 N$10723 N$10358 "Waveguide Crossing" sch_x=-58 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2689 N$10305 N$10307 N$10360 N$10362 "Waveguide Crossing" sch_x=-58 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2690 N$10309 N$10311 N$10364 N$10366 "Waveguide Crossing" sch_x=-58 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2691 N$10313 N$10315 N$10368 N$10370 "Waveguide Crossing" sch_x=-58 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2692 N$10317 N$10319 N$10372 N$10374 "Waveguide Crossing" sch_x=-58 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2693 N$10321 N$10323 N$10376 N$10378 "Waveguide Crossing" sch_x=-58 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2694 N$10325 N$10327 N$10380 N$10382 "Waveguide Crossing" sch_x=-58 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2695 N$10329 N$10331 N$10384 N$10386 "Waveguide Crossing" sch_x=-58 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2696 N$10333 N$10335 N$10388 N$10390 "Waveguide Crossing" sch_x=-58 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2697 N$10337 N$10339 N$10392 N$10394 "Waveguide Crossing" sch_x=-58 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2698 N$10341 N$10343 N$10396 N$10398 "Waveguide Crossing" sch_x=-58 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2699 N$10345 N$10347 N$10400 N$10402 "Waveguide Crossing" sch_x=-58 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2700 N$10349 N$10351 N$10404 N$10406 "Waveguide Crossing" sch_x=-58 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2701 N$10353 N$10355 N$10408 N$10777 "Waveguide Crossing" sch_x=-58 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2702 N$10357 N$10359 N$10725 N$10410 "Waveguide Crossing" sch_x=-56 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2703 N$10361 N$10363 N$10412 N$10414 "Waveguide Crossing" sch_x=-56 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2704 N$10365 N$10367 N$10416 N$10418 "Waveguide Crossing" sch_x=-56 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2705 N$10369 N$10371 N$10420 N$10422 "Waveguide Crossing" sch_x=-56 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2706 N$10373 N$10375 N$10424 N$10426 "Waveguide Crossing" sch_x=-56 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2707 N$10377 N$10379 N$10428 N$10430 "Waveguide Crossing" sch_x=-56 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2708 N$10381 N$10383 N$10432 N$10434 "Waveguide Crossing" sch_x=-56 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2709 N$10385 N$10387 N$10436 N$10438 "Waveguide Crossing" sch_x=-56 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2710 N$10389 N$10391 N$10440 N$10442 "Waveguide Crossing" sch_x=-56 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2711 N$10393 N$10395 N$10444 N$10446 "Waveguide Crossing" sch_x=-56 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2712 N$10397 N$10399 N$10448 N$10450 "Waveguide Crossing" sch_x=-56 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2713 N$10401 N$10403 N$10452 N$10454 "Waveguide Crossing" sch_x=-56 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2714 N$10405 N$10407 N$10456 N$10775 "Waveguide Crossing" sch_x=-56 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2715 N$10409 N$10411 N$10727 N$10458 "Waveguide Crossing" sch_x=-54 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2716 N$10413 N$10415 N$10460 N$10462 "Waveguide Crossing" sch_x=-54 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2717 N$10417 N$10419 N$10464 N$10466 "Waveguide Crossing" sch_x=-54 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2718 N$10421 N$10423 N$10468 N$10470 "Waveguide Crossing" sch_x=-54 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2719 N$10425 N$10427 N$10472 N$10474 "Waveguide Crossing" sch_x=-54 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2720 N$10429 N$10431 N$10476 N$10478 "Waveguide Crossing" sch_x=-54 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2721 N$10433 N$10435 N$10480 N$10482 "Waveguide Crossing" sch_x=-54 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2722 N$10437 N$10439 N$10484 N$10486 "Waveguide Crossing" sch_x=-54 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2723 N$10441 N$10443 N$10488 N$10490 "Waveguide Crossing" sch_x=-54 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2724 N$10445 N$10447 N$10492 N$10494 "Waveguide Crossing" sch_x=-54 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2725 N$10449 N$10451 N$10496 N$10498 "Waveguide Crossing" sch_x=-54 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2726 N$10453 N$10455 N$10500 N$10773 "Waveguide Crossing" sch_x=-54 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2727 N$10457 N$10459 N$10729 N$10502 "Waveguide Crossing" sch_x=-52 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2728 N$10461 N$10463 N$10504 N$10506 "Waveguide Crossing" sch_x=-52 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2729 N$10465 N$10467 N$10508 N$10510 "Waveguide Crossing" sch_x=-52 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2730 N$10469 N$10471 N$10512 N$10514 "Waveguide Crossing" sch_x=-52 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2731 N$10473 N$10475 N$10516 N$10518 "Waveguide Crossing" sch_x=-52 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2732 N$10477 N$10479 N$10520 N$10522 "Waveguide Crossing" sch_x=-52 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2733 N$10481 N$10483 N$10524 N$10526 "Waveguide Crossing" sch_x=-52 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2734 N$10485 N$10487 N$10528 N$10530 "Waveguide Crossing" sch_x=-52 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2735 N$10489 N$10491 N$10532 N$10534 "Waveguide Crossing" sch_x=-52 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2736 N$10493 N$10495 N$10536 N$10538 "Waveguide Crossing" sch_x=-52 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2737 N$10497 N$10499 N$10540 N$10771 "Waveguide Crossing" sch_x=-52 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2738 N$10501 N$10503 N$10731 N$10542 "Waveguide Crossing" sch_x=-50 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2739 N$10505 N$10507 N$10544 N$10546 "Waveguide Crossing" sch_x=-50 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2740 N$10509 N$10511 N$10548 N$10550 "Waveguide Crossing" sch_x=-50 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2741 N$10513 N$10515 N$10552 N$10554 "Waveguide Crossing" sch_x=-50 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2742 N$10517 N$10519 N$10556 N$10558 "Waveguide Crossing" sch_x=-50 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2743 N$10521 N$10523 N$10560 N$10562 "Waveguide Crossing" sch_x=-50 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2744 N$10525 N$10527 N$10564 N$10566 "Waveguide Crossing" sch_x=-50 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2745 N$10529 N$10531 N$10568 N$10570 "Waveguide Crossing" sch_x=-50 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2746 N$10533 N$10535 N$10572 N$10574 "Waveguide Crossing" sch_x=-50 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2747 N$10537 N$10539 N$10576 N$10769 "Waveguide Crossing" sch_x=-50 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2748 N$10541 N$10543 N$10733 N$10578 "Waveguide Crossing" sch_x=-48 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2749 N$10545 N$10547 N$10580 N$10582 "Waveguide Crossing" sch_x=-48 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2750 N$10549 N$10551 N$10584 N$10586 "Waveguide Crossing" sch_x=-48 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2751 N$10553 N$10555 N$10588 N$10590 "Waveguide Crossing" sch_x=-48 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2752 N$10557 N$10559 N$10592 N$10594 "Waveguide Crossing" sch_x=-48 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2753 N$10561 N$10563 N$10596 N$10598 "Waveguide Crossing" sch_x=-48 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2754 N$10565 N$10567 N$10600 N$10602 "Waveguide Crossing" sch_x=-48 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2755 N$10569 N$10571 N$10604 N$10606 "Waveguide Crossing" sch_x=-48 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2756 N$10573 N$10575 N$10608 N$10767 "Waveguide Crossing" sch_x=-48 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2757 N$10577 N$10579 N$10735 N$10610 "Waveguide Crossing" sch_x=-46 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2758 N$10581 N$10583 N$10612 N$10614 "Waveguide Crossing" sch_x=-46 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2759 N$10585 N$10587 N$10616 N$10618 "Waveguide Crossing" sch_x=-46 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2760 N$10589 N$10591 N$10620 N$10622 "Waveguide Crossing" sch_x=-46 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2761 N$10593 N$10595 N$10624 N$10626 "Waveguide Crossing" sch_x=-46 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2762 N$10597 N$10599 N$10628 N$10630 "Waveguide Crossing" sch_x=-46 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2763 N$10601 N$10603 N$10632 N$10634 "Waveguide Crossing" sch_x=-46 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2764 N$10605 N$10607 N$10636 N$10765 "Waveguide Crossing" sch_x=-46 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2765 N$10609 N$10611 N$10737 N$10638 "Waveguide Crossing" sch_x=-44 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2766 N$10613 N$10615 N$10640 N$10642 "Waveguide Crossing" sch_x=-44 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2767 N$10617 N$10619 N$10644 N$10646 "Waveguide Crossing" sch_x=-44 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2768 N$10621 N$10623 N$10648 N$10650 "Waveguide Crossing" sch_x=-44 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2769 N$10625 N$10627 N$10652 N$10654 "Waveguide Crossing" sch_x=-44 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2770 N$10629 N$10631 N$10656 N$10658 "Waveguide Crossing" sch_x=-44 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2771 N$10633 N$10635 N$10660 N$10763 "Waveguide Crossing" sch_x=-44 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2772 N$10637 N$10639 N$10739 N$10662 "Waveguide Crossing" sch_x=-42 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2773 N$10641 N$10643 N$10664 N$10666 "Waveguide Crossing" sch_x=-42 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2774 N$10645 N$10647 N$10668 N$10670 "Waveguide Crossing" sch_x=-42 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2775 N$10649 N$10651 N$10672 N$10674 "Waveguide Crossing" sch_x=-42 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2776 N$10653 N$10655 N$10676 N$10678 "Waveguide Crossing" sch_x=-42 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2777 N$10657 N$10659 N$10680 N$10761 "Waveguide Crossing" sch_x=-42 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2778 N$10661 N$10663 N$10741 N$10682 "Waveguide Crossing" sch_x=-40 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2779 N$10665 N$10667 N$10684 N$10686 "Waveguide Crossing" sch_x=-40 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2780 N$10669 N$10671 N$10688 N$10690 "Waveguide Crossing" sch_x=-40 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2781 N$10673 N$10675 N$10692 N$10694 "Waveguide Crossing" sch_x=-40 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2782 N$10677 N$10679 N$10696 N$10759 "Waveguide Crossing" sch_x=-40 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2783 N$10681 N$10683 N$10743 N$10698 "Waveguide Crossing" sch_x=-38 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2784 N$10685 N$10687 N$10700 N$10702 "Waveguide Crossing" sch_x=-38 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2785 N$10689 N$10691 N$10704 N$10706 "Waveguide Crossing" sch_x=-38 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2786 N$10693 N$10695 N$10708 N$10757 "Waveguide Crossing" sch_x=-38 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2787 N$10697 N$10699 N$10745 N$10710 "Waveguide Crossing" sch_x=-36 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2788 N$10701 N$10703 N$10712 N$10714 "Waveguide Crossing" sch_x=-36 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2789 N$10705 N$10707 N$10716 N$10755 "Waveguide Crossing" sch_x=-36 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2790 N$10709 N$10711 N$10747 N$10718 "Waveguide Crossing" sch_x=-34 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2791 N$10713 N$10715 N$10720 N$10753 "Waveguide Crossing" sch_x=-34 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2792 N$10717 N$10719 N$10749 N$10751 "Waveguide Crossing" sch_x=-32 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2585 N$10752 N$10754 N$10093 N$9954 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2586 N$10756 N$10758 N$9956 N$9958 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2587 N$10760 N$10762 N$9960 N$9962 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2588 N$10764 N$10766 N$9964 N$9966 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2589 N$10768 N$10770 N$9968 N$9970 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2590 N$10772 N$10774 N$9972 N$9974 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2591 N$10776 N$10778 N$9976 N$9978 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2592 N$10780 N$10784 N$9980 N$10095 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2593 N$9953 N$9955 N$10065 N$9982 "Waveguide Crossing" sch_x=-28 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2594 N$9957 N$9959 N$9984 N$9986 "Waveguide Crossing" sch_x=-28 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2595 N$9961 N$9963 N$9988 N$9990 "Waveguide Crossing" sch_x=-28 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2596 N$9965 N$9967 N$9992 N$9994 "Waveguide Crossing" sch_x=-28 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2597 N$9969 N$9971 N$9996 N$9998 "Waveguide Crossing" sch_x=-28 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2598 N$9973 N$9975 N$10000 N$10002 "Waveguide Crossing" sch_x=-28 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2599 N$9977 N$9979 N$10004 N$10091 "Waveguide Crossing" sch_x=-28 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2600 N$9981 N$9983 N$10067 N$10006 "Waveguide Crossing" sch_x=-26 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2601 N$9985 N$9987 N$10008 N$10010 "Waveguide Crossing" sch_x=-26 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2602 N$9989 N$9991 N$10012 N$10014 "Waveguide Crossing" sch_x=-26 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2603 N$9993 N$9995 N$10016 N$10018 "Waveguide Crossing" sch_x=-26 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2604 N$9997 N$9999 N$10020 N$10022 "Waveguide Crossing" sch_x=-26 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2605 N$10001 N$10003 N$10024 N$10089 "Waveguide Crossing" sch_x=-26 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2606 N$10005 N$10007 N$10069 N$10026 "Waveguide Crossing" sch_x=-24 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2607 N$10009 N$10011 N$10028 N$10030 "Waveguide Crossing" sch_x=-24 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2608 N$10013 N$10015 N$10032 N$10034 "Waveguide Crossing" sch_x=-24 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2609 N$10017 N$10019 N$10036 N$10038 "Waveguide Crossing" sch_x=-24 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2610 N$10021 N$10023 N$10040 N$10087 "Waveguide Crossing" sch_x=-24 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2611 N$10025 N$10027 N$10071 N$10042 "Waveguide Crossing" sch_x=-22 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2612 N$10029 N$10031 N$10044 N$10046 "Waveguide Crossing" sch_x=-22 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2613 N$10033 N$10035 N$10048 N$10050 "Waveguide Crossing" sch_x=-22 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2614 N$10037 N$10039 N$10052 N$10085 "Waveguide Crossing" sch_x=-22 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2615 N$10041 N$10043 N$10073 N$10054 "Waveguide Crossing" sch_x=-20 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2616 N$10045 N$10047 N$10056 N$10058 "Waveguide Crossing" sch_x=-20 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2617 N$10049 N$10051 N$10060 N$10083 "Waveguide Crossing" sch_x=-20 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2618 N$10053 N$10055 N$10075 N$10062 "Waveguide Crossing" sch_x=-18 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2619 N$10057 N$10059 N$10064 N$10081 "Waveguide Crossing" sch_x=-18 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2620 N$10061 N$10063 N$10077 N$10079 "Waveguide Crossing" sch_x=-16 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2565 N$10080 N$10082 N$9909 N$9874 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2566 N$10084 N$10086 N$9876 N$9878 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2567 N$10088 N$10090 N$9880 N$9882 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2568 N$10092 N$10096 N$9884 N$9911 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2569 N$9873 N$9875 N$9897 N$9886 "Waveguide Crossing" sch_x=-12 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2570 N$9877 N$9879 N$9888 N$9890 "Waveguide Crossing" sch_x=-12 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2571 N$9881 N$9883 N$9892 N$9907 "Waveguide Crossing" sch_x=-12 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2572 N$9885 N$9887 N$9899 N$9894 "Waveguide Crossing" sch_x=-10 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2573 N$9889 N$9891 N$9896 N$9905 "Waveguide Crossing" sch_x=-10 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2574 N$9893 N$9895 N$9901 N$9903 "Waveguide Crossing" sch_x=-8 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2513 N$10094 N$10066 N$9733 N$9698 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2514 N$10068 N$10070 N$9700 N$9702 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2515 N$10072 N$10074 N$9704 N$9706 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2516 N$10076 N$10078 N$9708 N$9735 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2517 N$9697 N$9699 N$9721 N$9710 "Waveguide Crossing" sch_x=-12 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2518 N$9701 N$9703 N$9712 N$9714 "Waveguide Crossing" sch_x=-12 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2519 N$9705 N$9707 N$9716 N$9731 "Waveguide Crossing" sch_x=-12 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2520 N$9709 N$9711 N$9723 N$9718 "Waveguide Crossing" sch_x=-10 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2521 N$9713 N$9715 N$9720 N$9729 "Waveguide Crossing" sch_x=-10 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2522 N$9717 N$9719 N$9725 N$9727 "Waveguide Crossing" sch_x=-8 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2409 N$10782 N$10722 N$9453 N$9314 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2410 N$10724 N$10726 N$9316 N$9318 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2411 N$10728 N$10730 N$9320 N$9322 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2412 N$10732 N$10734 N$9324 N$9326 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2413 N$10736 N$10738 N$9328 N$9330 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2414 N$10740 N$10742 N$9332 N$9334 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2415 N$10744 N$10746 N$9336 N$9338 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2416 N$10748 N$10750 N$9340 N$9455 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2417 N$9313 N$9315 N$9425 N$9342 "Waveguide Crossing" sch_x=-28 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2418 N$9317 N$9319 N$9344 N$9346 "Waveguide Crossing" sch_x=-28 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2419 N$9321 N$9323 N$9348 N$9350 "Waveguide Crossing" sch_x=-28 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2420 N$9325 N$9327 N$9352 N$9354 "Waveguide Crossing" sch_x=-28 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2421 N$9329 N$9331 N$9356 N$9358 "Waveguide Crossing" sch_x=-28 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2422 N$9333 N$9335 N$9360 N$9362 "Waveguide Crossing" sch_x=-28 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2423 N$9337 N$9339 N$9364 N$9451 "Waveguide Crossing" sch_x=-28 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2424 N$9341 N$9343 N$9427 N$9366 "Waveguide Crossing" sch_x=-26 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2425 N$9345 N$9347 N$9368 N$9370 "Waveguide Crossing" sch_x=-26 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2426 N$9349 N$9351 N$9372 N$9374 "Waveguide Crossing" sch_x=-26 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2427 N$9353 N$9355 N$9376 N$9378 "Waveguide Crossing" sch_x=-26 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2428 N$9357 N$9359 N$9380 N$9382 "Waveguide Crossing" sch_x=-26 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2429 N$9361 N$9363 N$9384 N$9449 "Waveguide Crossing" sch_x=-26 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2430 N$9365 N$9367 N$9429 N$9386 "Waveguide Crossing" sch_x=-24 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2431 N$9369 N$9371 N$9388 N$9390 "Waveguide Crossing" sch_x=-24 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2432 N$9373 N$9375 N$9392 N$9394 "Waveguide Crossing" sch_x=-24 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2433 N$9377 N$9379 N$9396 N$9398 "Waveguide Crossing" sch_x=-24 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2434 N$9381 N$9383 N$9400 N$9447 "Waveguide Crossing" sch_x=-24 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2435 N$9385 N$9387 N$9431 N$9402 "Waveguide Crossing" sch_x=-22 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2436 N$9389 N$9391 N$9404 N$9406 "Waveguide Crossing" sch_x=-22 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2437 N$9393 N$9395 N$9408 N$9410 "Waveguide Crossing" sch_x=-22 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2438 N$9397 N$9399 N$9412 N$9445 "Waveguide Crossing" sch_x=-22 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2439 N$9401 N$9403 N$9433 N$9414 "Waveguide Crossing" sch_x=-20 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2440 N$9405 N$9407 N$9416 N$9418 "Waveguide Crossing" sch_x=-20 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2441 N$9409 N$9411 N$9420 N$9443 "Waveguide Crossing" sch_x=-20 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2442 N$9413 N$9415 N$9435 N$9422 "Waveguide Crossing" sch_x=-18 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2443 N$9417 N$9419 N$9424 N$9441 "Waveguide Crossing" sch_x=-18 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2444 N$9421 N$9423 N$9437 N$9439 "Waveguide Crossing" sch_x=-16 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2389 N$9440 N$9442 N$9269 N$9234 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2390 N$9444 N$9446 N$9236 N$9238 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2391 N$9448 N$9450 N$9240 N$9242 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2392 N$9452 N$9456 N$9244 N$9271 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2393 N$9233 N$9235 N$9257 N$9246 "Waveguide Crossing" sch_x=-12 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2394 N$9237 N$9239 N$9248 N$9250 "Waveguide Crossing" sch_x=-12 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2395 N$9241 N$9243 N$9252 N$9267 "Waveguide Crossing" sch_x=-12 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2396 N$9245 N$9247 N$9259 N$9254 "Waveguide Crossing" sch_x=-10 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2397 N$9249 N$9251 N$9256 N$9265 "Waveguide Crossing" sch_x=-10 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2398 N$9253 N$9255 N$9261 N$9263 "Waveguide Crossing" sch_x=-8 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2337 N$9454 N$9426 N$9093 N$9058 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2338 N$9428 N$9430 N$9060 N$9062 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2339 N$9432 N$9434 N$9064 N$9066 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2340 N$9436 N$9438 N$9068 N$9095 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2341 N$9057 N$9059 N$9081 N$9070 "Waveguide Crossing" sch_x=-12 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2342 N$9061 N$9063 N$9072 N$9074 "Waveguide Crossing" sch_x=-12 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2343 N$9065 N$9067 N$9076 N$9091 "Waveguide Crossing" sch_x=-12 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2344 N$9069 N$9071 N$9083 N$9078 "Waveguide Crossing" sch_x=-10 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2345 N$9073 N$9075 N$9080 N$9089 "Waveguide Crossing" sch_x=-10 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2346 N$9077 N$9079 N$9085 N$9087 "Waveguide Crossing" sch_x=-8 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1249 N$26238 N$25986 N$6845 N$4738 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1250 N$25988 N$25990 N$4740 N$4742 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1251 N$25992 N$25994 N$4744 N$4746 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1252 N$25996 N$25998 N$4748 N$4750 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1253 N$26000 N$26002 N$4752 N$4754 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1254 N$26004 N$26006 N$4756 N$4758 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1255 N$26008 N$26010 N$4760 N$4762 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1256 N$26012 N$26014 N$4764 N$4766 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1257 N$26016 N$26018 N$4768 N$4770 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1258 N$26020 N$26022 N$4772 N$4774 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1259 N$26024 N$26026 N$4776 N$4778 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1260 N$26028 N$26030 N$4780 N$4782 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1261 N$26032 N$26034 N$4784 N$4786 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1262 N$26036 N$26038 N$4788 N$4790 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1263 N$26040 N$26042 N$4792 N$4794 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1264 N$26044 N$26046 N$4796 N$4798 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1265 N$26048 N$26050 N$4800 N$4802 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1266 N$26052 N$26054 N$4804 N$4806 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1267 N$26056 N$26058 N$4808 N$4810 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1268 N$26060 N$26062 N$4812 N$4814 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1269 N$26064 N$26066 N$4816 N$4818 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1270 N$26068 N$26070 N$4820 N$4822 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1271 N$26072 N$26074 N$4824 N$4826 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1272 N$26076 N$26078 N$4828 N$4830 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1273 N$26080 N$26082 N$4832 N$4834 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1274 N$26084 N$26086 N$4836 N$4838 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1275 N$26088 N$26090 N$4840 N$4842 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1276 N$26092 N$26094 N$4844 N$4846 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1277 N$26096 N$26098 N$4848 N$4850 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1278 N$26100 N$26102 N$4852 N$4854 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1279 N$26104 N$26106 N$4856 N$4858 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1280 N$26108 N$26110 N$4860 N$6847 BDC_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1281 N$4737 N$4739 N$6721 N$4862 "Waveguide Crossing" sch_x=-124 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1282 N$4741 N$4743 N$4864 N$4866 "Waveguide Crossing" sch_x=-124 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1283 N$4745 N$4747 N$4868 N$4870 "Waveguide Crossing" sch_x=-124 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1284 N$4749 N$4751 N$4872 N$4874 "Waveguide Crossing" sch_x=-124 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1285 N$4753 N$4755 N$4876 N$4878 "Waveguide Crossing" sch_x=-124 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1286 N$4757 N$4759 N$4880 N$4882 "Waveguide Crossing" sch_x=-124 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1287 N$4761 N$4763 N$4884 N$4886 "Waveguide Crossing" sch_x=-124 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1288 N$4765 N$4767 N$4888 N$4890 "Waveguide Crossing" sch_x=-124 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1289 N$4769 N$4771 N$4892 N$4894 "Waveguide Crossing" sch_x=-124 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1290 N$4773 N$4775 N$4896 N$4898 "Waveguide Crossing" sch_x=-124 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1291 N$4777 N$4779 N$4900 N$4902 "Waveguide Crossing" sch_x=-124 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1292 N$4781 N$4783 N$4904 N$4906 "Waveguide Crossing" sch_x=-124 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1293 N$4785 N$4787 N$4908 N$4910 "Waveguide Crossing" sch_x=-124 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1294 N$4789 N$4791 N$4912 N$4914 "Waveguide Crossing" sch_x=-124 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1295 N$4793 N$4795 N$4916 N$4918 "Waveguide Crossing" sch_x=-124 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1296 N$4797 N$4799 N$4920 N$4922 "Waveguide Crossing" sch_x=-124 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1297 N$4801 N$4803 N$4924 N$4926 "Waveguide Crossing" sch_x=-124 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1298 N$4805 N$4807 N$4928 N$4930 "Waveguide Crossing" sch_x=-124 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1299 N$4809 N$4811 N$4932 N$4934 "Waveguide Crossing" sch_x=-124 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1300 N$4813 N$4815 N$4936 N$4938 "Waveguide Crossing" sch_x=-124 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1301 N$4817 N$4819 N$4940 N$4942 "Waveguide Crossing" sch_x=-124 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1302 N$4821 N$4823 N$4944 N$4946 "Waveguide Crossing" sch_x=-124 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1303 N$4825 N$4827 N$4948 N$4950 "Waveguide Crossing" sch_x=-124 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1304 N$4829 N$4831 N$4952 N$4954 "Waveguide Crossing" sch_x=-124 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1305 N$4833 N$4835 N$4956 N$4958 "Waveguide Crossing" sch_x=-124 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1306 N$4837 N$4839 N$4960 N$4962 "Waveguide Crossing" sch_x=-124 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1307 N$4841 N$4843 N$4964 N$4966 "Waveguide Crossing" sch_x=-124 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1308 N$4845 N$4847 N$4968 N$4970 "Waveguide Crossing" sch_x=-124 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1309 N$4849 N$4851 N$4972 N$4974 "Waveguide Crossing" sch_x=-124 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1310 N$4853 N$4855 N$4976 N$4978 "Waveguide Crossing" sch_x=-124 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1311 N$4857 N$4859 N$4980 N$6843 "Waveguide Crossing" sch_x=-124 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1312 N$4861 N$4863 N$6723 N$4982 "Waveguide Crossing" sch_x=-122 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1313 N$4865 N$4867 N$4984 N$4986 "Waveguide Crossing" sch_x=-122 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1314 N$4869 N$4871 N$4988 N$4990 "Waveguide Crossing" sch_x=-122 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1315 N$4873 N$4875 N$4992 N$4994 "Waveguide Crossing" sch_x=-122 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1316 N$4877 N$4879 N$4996 N$4998 "Waveguide Crossing" sch_x=-122 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1317 N$4881 N$4883 N$5000 N$5002 "Waveguide Crossing" sch_x=-122 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1318 N$4885 N$4887 N$5004 N$5006 "Waveguide Crossing" sch_x=-122 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1319 N$4889 N$4891 N$5008 N$5010 "Waveguide Crossing" sch_x=-122 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1320 N$4893 N$4895 N$5012 N$5014 "Waveguide Crossing" sch_x=-122 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1321 N$4897 N$4899 N$5016 N$5018 "Waveguide Crossing" sch_x=-122 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1322 N$4901 N$4903 N$5020 N$5022 "Waveguide Crossing" sch_x=-122 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1323 N$4905 N$4907 N$5024 N$5026 "Waveguide Crossing" sch_x=-122 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1324 N$4909 N$4911 N$5028 N$5030 "Waveguide Crossing" sch_x=-122 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1325 N$4913 N$4915 N$5032 N$5034 "Waveguide Crossing" sch_x=-122 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1326 N$4917 N$4919 N$5036 N$5038 "Waveguide Crossing" sch_x=-122 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1327 N$4921 N$4923 N$5040 N$5042 "Waveguide Crossing" sch_x=-122 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1328 N$4925 N$4927 N$5044 N$5046 "Waveguide Crossing" sch_x=-122 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1329 N$4929 N$4931 N$5048 N$5050 "Waveguide Crossing" sch_x=-122 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1330 N$4933 N$4935 N$5052 N$5054 "Waveguide Crossing" sch_x=-122 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1331 N$4937 N$4939 N$5056 N$5058 "Waveguide Crossing" sch_x=-122 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1332 N$4941 N$4943 N$5060 N$5062 "Waveguide Crossing" sch_x=-122 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1333 N$4945 N$4947 N$5064 N$5066 "Waveguide Crossing" sch_x=-122 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1334 N$4949 N$4951 N$5068 N$5070 "Waveguide Crossing" sch_x=-122 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1335 N$4953 N$4955 N$5072 N$5074 "Waveguide Crossing" sch_x=-122 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1336 N$4957 N$4959 N$5076 N$5078 "Waveguide Crossing" sch_x=-122 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1337 N$4961 N$4963 N$5080 N$5082 "Waveguide Crossing" sch_x=-122 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1338 N$4965 N$4967 N$5084 N$5086 "Waveguide Crossing" sch_x=-122 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1339 N$4969 N$4971 N$5088 N$5090 "Waveguide Crossing" sch_x=-122 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1340 N$4973 N$4975 N$5092 N$5094 "Waveguide Crossing" sch_x=-122 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1341 N$4977 N$4979 N$5096 N$6841 "Waveguide Crossing" sch_x=-122 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1342 N$4981 N$4983 N$6725 N$5098 "Waveguide Crossing" sch_x=-120 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1343 N$4985 N$4987 N$5100 N$5102 "Waveguide Crossing" sch_x=-120 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1344 N$4989 N$4991 N$5104 N$5106 "Waveguide Crossing" sch_x=-120 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1345 N$4993 N$4995 N$5108 N$5110 "Waveguide Crossing" sch_x=-120 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1346 N$4997 N$4999 N$5112 N$5114 "Waveguide Crossing" sch_x=-120 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1347 N$5001 N$5003 N$5116 N$5118 "Waveguide Crossing" sch_x=-120 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1348 N$5005 N$5007 N$5120 N$5122 "Waveguide Crossing" sch_x=-120 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1349 N$5009 N$5011 N$5124 N$5126 "Waveguide Crossing" sch_x=-120 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1350 N$5013 N$5015 N$5128 N$5130 "Waveguide Crossing" sch_x=-120 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1351 N$5017 N$5019 N$5132 N$5134 "Waveguide Crossing" sch_x=-120 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1352 N$5021 N$5023 N$5136 N$5138 "Waveguide Crossing" sch_x=-120 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1353 N$5025 N$5027 N$5140 N$5142 "Waveguide Crossing" sch_x=-120 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1354 N$5029 N$5031 N$5144 N$5146 "Waveguide Crossing" sch_x=-120 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1355 N$5033 N$5035 N$5148 N$5150 "Waveguide Crossing" sch_x=-120 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1356 N$5037 N$5039 N$5152 N$5154 "Waveguide Crossing" sch_x=-120 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1357 N$5041 N$5043 N$5156 N$5158 "Waveguide Crossing" sch_x=-120 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1358 N$5045 N$5047 N$5160 N$5162 "Waveguide Crossing" sch_x=-120 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1359 N$5049 N$5051 N$5164 N$5166 "Waveguide Crossing" sch_x=-120 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1360 N$5053 N$5055 N$5168 N$5170 "Waveguide Crossing" sch_x=-120 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1361 N$5057 N$5059 N$5172 N$5174 "Waveguide Crossing" sch_x=-120 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1362 N$5061 N$5063 N$5176 N$5178 "Waveguide Crossing" sch_x=-120 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1363 N$5065 N$5067 N$5180 N$5182 "Waveguide Crossing" sch_x=-120 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1364 N$5069 N$5071 N$5184 N$5186 "Waveguide Crossing" sch_x=-120 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1365 N$5073 N$5075 N$5188 N$5190 "Waveguide Crossing" sch_x=-120 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1366 N$5077 N$5079 N$5192 N$5194 "Waveguide Crossing" sch_x=-120 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1367 N$5081 N$5083 N$5196 N$5198 "Waveguide Crossing" sch_x=-120 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1368 N$5085 N$5087 N$5200 N$5202 "Waveguide Crossing" sch_x=-120 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1369 N$5089 N$5091 N$5204 N$5206 "Waveguide Crossing" sch_x=-120 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1370 N$5093 N$5095 N$5208 N$6839 "Waveguide Crossing" sch_x=-120 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1371 N$5097 N$5099 N$6727 N$5210 "Waveguide Crossing" sch_x=-118 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1372 N$5101 N$5103 N$5212 N$5214 "Waveguide Crossing" sch_x=-118 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1373 N$5105 N$5107 N$5216 N$5218 "Waveguide Crossing" sch_x=-118 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1374 N$5109 N$5111 N$5220 N$5222 "Waveguide Crossing" sch_x=-118 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1375 N$5113 N$5115 N$5224 N$5226 "Waveguide Crossing" sch_x=-118 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1376 N$5117 N$5119 N$5228 N$5230 "Waveguide Crossing" sch_x=-118 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1377 N$5121 N$5123 N$5232 N$5234 "Waveguide Crossing" sch_x=-118 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1378 N$5125 N$5127 N$5236 N$5238 "Waveguide Crossing" sch_x=-118 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1379 N$5129 N$5131 N$5240 N$5242 "Waveguide Crossing" sch_x=-118 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1380 N$5133 N$5135 N$5244 N$5246 "Waveguide Crossing" sch_x=-118 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1381 N$5137 N$5139 N$5248 N$5250 "Waveguide Crossing" sch_x=-118 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1382 N$5141 N$5143 N$5252 N$5254 "Waveguide Crossing" sch_x=-118 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1383 N$5145 N$5147 N$5256 N$5258 "Waveguide Crossing" sch_x=-118 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1384 N$5149 N$5151 N$5260 N$5262 "Waveguide Crossing" sch_x=-118 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1385 N$5153 N$5155 N$5264 N$5266 "Waveguide Crossing" sch_x=-118 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1386 N$5157 N$5159 N$5268 N$5270 "Waveguide Crossing" sch_x=-118 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1387 N$5161 N$5163 N$5272 N$5274 "Waveguide Crossing" sch_x=-118 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1388 N$5165 N$5167 N$5276 N$5278 "Waveguide Crossing" sch_x=-118 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1389 N$5169 N$5171 N$5280 N$5282 "Waveguide Crossing" sch_x=-118 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1390 N$5173 N$5175 N$5284 N$5286 "Waveguide Crossing" sch_x=-118 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1391 N$5177 N$5179 N$5288 N$5290 "Waveguide Crossing" sch_x=-118 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1392 N$5181 N$5183 N$5292 N$5294 "Waveguide Crossing" sch_x=-118 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1393 N$5185 N$5187 N$5296 N$5298 "Waveguide Crossing" sch_x=-118 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1394 N$5189 N$5191 N$5300 N$5302 "Waveguide Crossing" sch_x=-118 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1395 N$5193 N$5195 N$5304 N$5306 "Waveguide Crossing" sch_x=-118 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1396 N$5197 N$5199 N$5308 N$5310 "Waveguide Crossing" sch_x=-118 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1397 N$5201 N$5203 N$5312 N$5314 "Waveguide Crossing" sch_x=-118 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1398 N$5205 N$5207 N$5316 N$6837 "Waveguide Crossing" sch_x=-118 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1399 N$5209 N$5211 N$6729 N$5318 "Waveguide Crossing" sch_x=-116 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1400 N$5213 N$5215 N$5320 N$5322 "Waveguide Crossing" sch_x=-116 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1401 N$5217 N$5219 N$5324 N$5326 "Waveguide Crossing" sch_x=-116 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1402 N$5221 N$5223 N$5328 N$5330 "Waveguide Crossing" sch_x=-116 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1403 N$5225 N$5227 N$5332 N$5334 "Waveguide Crossing" sch_x=-116 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1404 N$5229 N$5231 N$5336 N$5338 "Waveguide Crossing" sch_x=-116 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1405 N$5233 N$5235 N$5340 N$5342 "Waveguide Crossing" sch_x=-116 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1406 N$5237 N$5239 N$5344 N$5346 "Waveguide Crossing" sch_x=-116 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1407 N$5241 N$5243 N$5348 N$5350 "Waveguide Crossing" sch_x=-116 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1408 N$5245 N$5247 N$5352 N$5354 "Waveguide Crossing" sch_x=-116 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1409 N$5249 N$5251 N$5356 N$5358 "Waveguide Crossing" sch_x=-116 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1410 N$5253 N$5255 N$5360 N$5362 "Waveguide Crossing" sch_x=-116 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1411 N$5257 N$5259 N$5364 N$5366 "Waveguide Crossing" sch_x=-116 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1412 N$5261 N$5263 N$5368 N$5370 "Waveguide Crossing" sch_x=-116 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1413 N$5265 N$5267 N$5372 N$5374 "Waveguide Crossing" sch_x=-116 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1414 N$5269 N$5271 N$5376 N$5378 "Waveguide Crossing" sch_x=-116 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1415 N$5273 N$5275 N$5380 N$5382 "Waveguide Crossing" sch_x=-116 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1416 N$5277 N$5279 N$5384 N$5386 "Waveguide Crossing" sch_x=-116 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1417 N$5281 N$5283 N$5388 N$5390 "Waveguide Crossing" sch_x=-116 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1418 N$5285 N$5287 N$5392 N$5394 "Waveguide Crossing" sch_x=-116 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1419 N$5289 N$5291 N$5396 N$5398 "Waveguide Crossing" sch_x=-116 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1420 N$5293 N$5295 N$5400 N$5402 "Waveguide Crossing" sch_x=-116 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1421 N$5297 N$5299 N$5404 N$5406 "Waveguide Crossing" sch_x=-116 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1422 N$5301 N$5303 N$5408 N$5410 "Waveguide Crossing" sch_x=-116 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1423 N$5305 N$5307 N$5412 N$5414 "Waveguide Crossing" sch_x=-116 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1424 N$5309 N$5311 N$5416 N$5418 "Waveguide Crossing" sch_x=-116 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1425 N$5313 N$5315 N$5420 N$6835 "Waveguide Crossing" sch_x=-116 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1426 N$5317 N$5319 N$6731 N$5422 "Waveguide Crossing" sch_x=-114 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1427 N$5321 N$5323 N$5424 N$5426 "Waveguide Crossing" sch_x=-114 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1428 N$5325 N$5327 N$5428 N$5430 "Waveguide Crossing" sch_x=-114 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1429 N$5329 N$5331 N$5432 N$5434 "Waveguide Crossing" sch_x=-114 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1430 N$5333 N$5335 N$5436 N$5438 "Waveguide Crossing" sch_x=-114 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1431 N$5337 N$5339 N$5440 N$5442 "Waveguide Crossing" sch_x=-114 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1432 N$5341 N$5343 N$5444 N$5446 "Waveguide Crossing" sch_x=-114 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1433 N$5345 N$5347 N$5448 N$5450 "Waveguide Crossing" sch_x=-114 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1434 N$5349 N$5351 N$5452 N$5454 "Waveguide Crossing" sch_x=-114 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1435 N$5353 N$5355 N$5456 N$5458 "Waveguide Crossing" sch_x=-114 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1436 N$5357 N$5359 N$5460 N$5462 "Waveguide Crossing" sch_x=-114 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1437 N$5361 N$5363 N$5464 N$5466 "Waveguide Crossing" sch_x=-114 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1438 N$5365 N$5367 N$5468 N$5470 "Waveguide Crossing" sch_x=-114 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1439 N$5369 N$5371 N$5472 N$5474 "Waveguide Crossing" sch_x=-114 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1440 N$5373 N$5375 N$5476 N$5478 "Waveguide Crossing" sch_x=-114 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1441 N$5377 N$5379 N$5480 N$5482 "Waveguide Crossing" sch_x=-114 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1442 N$5381 N$5383 N$5484 N$5486 "Waveguide Crossing" sch_x=-114 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1443 N$5385 N$5387 N$5488 N$5490 "Waveguide Crossing" sch_x=-114 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1444 N$5389 N$5391 N$5492 N$5494 "Waveguide Crossing" sch_x=-114 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1445 N$5393 N$5395 N$5496 N$5498 "Waveguide Crossing" sch_x=-114 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1446 N$5397 N$5399 N$5500 N$5502 "Waveguide Crossing" sch_x=-114 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1447 N$5401 N$5403 N$5504 N$5506 "Waveguide Crossing" sch_x=-114 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1448 N$5405 N$5407 N$5508 N$5510 "Waveguide Crossing" sch_x=-114 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1449 N$5409 N$5411 N$5512 N$5514 "Waveguide Crossing" sch_x=-114 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1450 N$5413 N$5415 N$5516 N$5518 "Waveguide Crossing" sch_x=-114 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1451 N$5417 N$5419 N$5520 N$6833 "Waveguide Crossing" sch_x=-114 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1452 N$5421 N$5423 N$6733 N$5522 "Waveguide Crossing" sch_x=-112 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1453 N$5425 N$5427 N$5524 N$5526 "Waveguide Crossing" sch_x=-112 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1454 N$5429 N$5431 N$5528 N$5530 "Waveguide Crossing" sch_x=-112 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1455 N$5433 N$5435 N$5532 N$5534 "Waveguide Crossing" sch_x=-112 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1456 N$5437 N$5439 N$5536 N$5538 "Waveguide Crossing" sch_x=-112 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1457 N$5441 N$5443 N$5540 N$5542 "Waveguide Crossing" sch_x=-112 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1458 N$5445 N$5447 N$5544 N$5546 "Waveguide Crossing" sch_x=-112 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1459 N$5449 N$5451 N$5548 N$5550 "Waveguide Crossing" sch_x=-112 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1460 N$5453 N$5455 N$5552 N$5554 "Waveguide Crossing" sch_x=-112 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1461 N$5457 N$5459 N$5556 N$5558 "Waveguide Crossing" sch_x=-112 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1462 N$5461 N$5463 N$5560 N$5562 "Waveguide Crossing" sch_x=-112 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1463 N$5465 N$5467 N$5564 N$5566 "Waveguide Crossing" sch_x=-112 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1464 N$5469 N$5471 N$5568 N$5570 "Waveguide Crossing" sch_x=-112 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1465 N$5473 N$5475 N$5572 N$5574 "Waveguide Crossing" sch_x=-112 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1466 N$5477 N$5479 N$5576 N$5578 "Waveguide Crossing" sch_x=-112 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1467 N$5481 N$5483 N$5580 N$5582 "Waveguide Crossing" sch_x=-112 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1468 N$5485 N$5487 N$5584 N$5586 "Waveguide Crossing" sch_x=-112 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1469 N$5489 N$5491 N$5588 N$5590 "Waveguide Crossing" sch_x=-112 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1470 N$5493 N$5495 N$5592 N$5594 "Waveguide Crossing" sch_x=-112 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1471 N$5497 N$5499 N$5596 N$5598 "Waveguide Crossing" sch_x=-112 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1472 N$5501 N$5503 N$5600 N$5602 "Waveguide Crossing" sch_x=-112 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1473 N$5505 N$5507 N$5604 N$5606 "Waveguide Crossing" sch_x=-112 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1474 N$5509 N$5511 N$5608 N$5610 "Waveguide Crossing" sch_x=-112 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1475 N$5513 N$5515 N$5612 N$5614 "Waveguide Crossing" sch_x=-112 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1476 N$5517 N$5519 N$5616 N$6831 "Waveguide Crossing" sch_x=-112 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1477 N$5521 N$5523 N$6735 N$5618 "Waveguide Crossing" sch_x=-110 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1478 N$5525 N$5527 N$5620 N$5622 "Waveguide Crossing" sch_x=-110 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1479 N$5529 N$5531 N$5624 N$5626 "Waveguide Crossing" sch_x=-110 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1480 N$5533 N$5535 N$5628 N$5630 "Waveguide Crossing" sch_x=-110 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1481 N$5537 N$5539 N$5632 N$5634 "Waveguide Crossing" sch_x=-110 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1482 N$5541 N$5543 N$5636 N$5638 "Waveguide Crossing" sch_x=-110 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1483 N$5545 N$5547 N$5640 N$5642 "Waveguide Crossing" sch_x=-110 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1484 N$5549 N$5551 N$5644 N$5646 "Waveguide Crossing" sch_x=-110 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1485 N$5553 N$5555 N$5648 N$5650 "Waveguide Crossing" sch_x=-110 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1486 N$5557 N$5559 N$5652 N$5654 "Waveguide Crossing" sch_x=-110 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1487 N$5561 N$5563 N$5656 N$5658 "Waveguide Crossing" sch_x=-110 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1488 N$5565 N$5567 N$5660 N$5662 "Waveguide Crossing" sch_x=-110 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1489 N$5569 N$5571 N$5664 N$5666 "Waveguide Crossing" sch_x=-110 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1490 N$5573 N$5575 N$5668 N$5670 "Waveguide Crossing" sch_x=-110 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1491 N$5577 N$5579 N$5672 N$5674 "Waveguide Crossing" sch_x=-110 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1492 N$5581 N$5583 N$5676 N$5678 "Waveguide Crossing" sch_x=-110 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1493 N$5585 N$5587 N$5680 N$5682 "Waveguide Crossing" sch_x=-110 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1494 N$5589 N$5591 N$5684 N$5686 "Waveguide Crossing" sch_x=-110 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1495 N$5593 N$5595 N$5688 N$5690 "Waveguide Crossing" sch_x=-110 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1496 N$5597 N$5599 N$5692 N$5694 "Waveguide Crossing" sch_x=-110 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1497 N$5601 N$5603 N$5696 N$5698 "Waveguide Crossing" sch_x=-110 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1498 N$5605 N$5607 N$5700 N$5702 "Waveguide Crossing" sch_x=-110 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1499 N$5609 N$5611 N$5704 N$5706 "Waveguide Crossing" sch_x=-110 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1500 N$5613 N$5615 N$5708 N$6829 "Waveguide Crossing" sch_x=-110 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1501 N$5617 N$5619 N$6737 N$5710 "Waveguide Crossing" sch_x=-108 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1502 N$5621 N$5623 N$5712 N$5714 "Waveguide Crossing" sch_x=-108 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1503 N$5625 N$5627 N$5716 N$5718 "Waveguide Crossing" sch_x=-108 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1504 N$5629 N$5631 N$5720 N$5722 "Waveguide Crossing" sch_x=-108 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1505 N$5633 N$5635 N$5724 N$5726 "Waveguide Crossing" sch_x=-108 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1506 N$5637 N$5639 N$5728 N$5730 "Waveguide Crossing" sch_x=-108 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1507 N$5641 N$5643 N$5732 N$5734 "Waveguide Crossing" sch_x=-108 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1508 N$5645 N$5647 N$5736 N$5738 "Waveguide Crossing" sch_x=-108 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1509 N$5649 N$5651 N$5740 N$5742 "Waveguide Crossing" sch_x=-108 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1510 N$5653 N$5655 N$5744 N$5746 "Waveguide Crossing" sch_x=-108 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1511 N$5657 N$5659 N$5748 N$5750 "Waveguide Crossing" sch_x=-108 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1512 N$5661 N$5663 N$5752 N$5754 "Waveguide Crossing" sch_x=-108 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1513 N$5665 N$5667 N$5756 N$5758 "Waveguide Crossing" sch_x=-108 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1514 N$5669 N$5671 N$5760 N$5762 "Waveguide Crossing" sch_x=-108 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1515 N$5673 N$5675 N$5764 N$5766 "Waveguide Crossing" sch_x=-108 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1516 N$5677 N$5679 N$5768 N$5770 "Waveguide Crossing" sch_x=-108 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1517 N$5681 N$5683 N$5772 N$5774 "Waveguide Crossing" sch_x=-108 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1518 N$5685 N$5687 N$5776 N$5778 "Waveguide Crossing" sch_x=-108 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1519 N$5689 N$5691 N$5780 N$5782 "Waveguide Crossing" sch_x=-108 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1520 N$5693 N$5695 N$5784 N$5786 "Waveguide Crossing" sch_x=-108 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1521 N$5697 N$5699 N$5788 N$5790 "Waveguide Crossing" sch_x=-108 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1522 N$5701 N$5703 N$5792 N$5794 "Waveguide Crossing" sch_x=-108 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1523 N$5705 N$5707 N$5796 N$6827 "Waveguide Crossing" sch_x=-108 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1524 N$5709 N$5711 N$6739 N$5798 "Waveguide Crossing" sch_x=-106 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1525 N$5713 N$5715 N$5800 N$5802 "Waveguide Crossing" sch_x=-106 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1526 N$5717 N$5719 N$5804 N$5806 "Waveguide Crossing" sch_x=-106 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1527 N$5721 N$5723 N$5808 N$5810 "Waveguide Crossing" sch_x=-106 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1528 N$5725 N$5727 N$5812 N$5814 "Waveguide Crossing" sch_x=-106 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1529 N$5729 N$5731 N$5816 N$5818 "Waveguide Crossing" sch_x=-106 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1530 N$5733 N$5735 N$5820 N$5822 "Waveguide Crossing" sch_x=-106 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1531 N$5737 N$5739 N$5824 N$5826 "Waveguide Crossing" sch_x=-106 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1532 N$5741 N$5743 N$5828 N$5830 "Waveguide Crossing" sch_x=-106 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1533 N$5745 N$5747 N$5832 N$5834 "Waveguide Crossing" sch_x=-106 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1534 N$5749 N$5751 N$5836 N$5838 "Waveguide Crossing" sch_x=-106 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1535 N$5753 N$5755 N$5840 N$5842 "Waveguide Crossing" sch_x=-106 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1536 N$5757 N$5759 N$5844 N$5846 "Waveguide Crossing" sch_x=-106 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1537 N$5761 N$5763 N$5848 N$5850 "Waveguide Crossing" sch_x=-106 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1538 N$5765 N$5767 N$5852 N$5854 "Waveguide Crossing" sch_x=-106 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1539 N$5769 N$5771 N$5856 N$5858 "Waveguide Crossing" sch_x=-106 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1540 N$5773 N$5775 N$5860 N$5862 "Waveguide Crossing" sch_x=-106 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1541 N$5777 N$5779 N$5864 N$5866 "Waveguide Crossing" sch_x=-106 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1542 N$5781 N$5783 N$5868 N$5870 "Waveguide Crossing" sch_x=-106 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1543 N$5785 N$5787 N$5872 N$5874 "Waveguide Crossing" sch_x=-106 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1544 N$5789 N$5791 N$5876 N$5878 "Waveguide Crossing" sch_x=-106 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1545 N$5793 N$5795 N$5880 N$6825 "Waveguide Crossing" sch_x=-106 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1546 N$5797 N$5799 N$6741 N$5882 "Waveguide Crossing" sch_x=-104 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1547 N$5801 N$5803 N$5884 N$5886 "Waveguide Crossing" sch_x=-104 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1548 N$5805 N$5807 N$5888 N$5890 "Waveguide Crossing" sch_x=-104 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1549 N$5809 N$5811 N$5892 N$5894 "Waveguide Crossing" sch_x=-104 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1550 N$5813 N$5815 N$5896 N$5898 "Waveguide Crossing" sch_x=-104 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1551 N$5817 N$5819 N$5900 N$5902 "Waveguide Crossing" sch_x=-104 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1552 N$5821 N$5823 N$5904 N$5906 "Waveguide Crossing" sch_x=-104 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1553 N$5825 N$5827 N$5908 N$5910 "Waveguide Crossing" sch_x=-104 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1554 N$5829 N$5831 N$5912 N$5914 "Waveguide Crossing" sch_x=-104 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1555 N$5833 N$5835 N$5916 N$5918 "Waveguide Crossing" sch_x=-104 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1556 N$5837 N$5839 N$5920 N$5922 "Waveguide Crossing" sch_x=-104 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1557 N$5841 N$5843 N$5924 N$5926 "Waveguide Crossing" sch_x=-104 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1558 N$5845 N$5847 N$5928 N$5930 "Waveguide Crossing" sch_x=-104 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1559 N$5849 N$5851 N$5932 N$5934 "Waveguide Crossing" sch_x=-104 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1560 N$5853 N$5855 N$5936 N$5938 "Waveguide Crossing" sch_x=-104 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1561 N$5857 N$5859 N$5940 N$5942 "Waveguide Crossing" sch_x=-104 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1562 N$5861 N$5863 N$5944 N$5946 "Waveguide Crossing" sch_x=-104 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1563 N$5865 N$5867 N$5948 N$5950 "Waveguide Crossing" sch_x=-104 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1564 N$5869 N$5871 N$5952 N$5954 "Waveguide Crossing" sch_x=-104 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1565 N$5873 N$5875 N$5956 N$5958 "Waveguide Crossing" sch_x=-104 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1566 N$5877 N$5879 N$5960 N$6823 "Waveguide Crossing" sch_x=-104 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1567 N$5881 N$5883 N$6743 N$5962 "Waveguide Crossing" sch_x=-102 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1568 N$5885 N$5887 N$5964 N$5966 "Waveguide Crossing" sch_x=-102 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1569 N$5889 N$5891 N$5968 N$5970 "Waveguide Crossing" sch_x=-102 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1570 N$5893 N$5895 N$5972 N$5974 "Waveguide Crossing" sch_x=-102 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1571 N$5897 N$5899 N$5976 N$5978 "Waveguide Crossing" sch_x=-102 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1572 N$5901 N$5903 N$5980 N$5982 "Waveguide Crossing" sch_x=-102 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1573 N$5905 N$5907 N$5984 N$5986 "Waveguide Crossing" sch_x=-102 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1574 N$5909 N$5911 N$5988 N$5990 "Waveguide Crossing" sch_x=-102 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1575 N$5913 N$5915 N$5992 N$5994 "Waveguide Crossing" sch_x=-102 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1576 N$5917 N$5919 N$5996 N$5998 "Waveguide Crossing" sch_x=-102 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1577 N$5921 N$5923 N$6000 N$6002 "Waveguide Crossing" sch_x=-102 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1578 N$5925 N$5927 N$6004 N$6006 "Waveguide Crossing" sch_x=-102 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1579 N$5929 N$5931 N$6008 N$6010 "Waveguide Crossing" sch_x=-102 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1580 N$5933 N$5935 N$6012 N$6014 "Waveguide Crossing" sch_x=-102 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1581 N$5937 N$5939 N$6016 N$6018 "Waveguide Crossing" sch_x=-102 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1582 N$5941 N$5943 N$6020 N$6022 "Waveguide Crossing" sch_x=-102 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1583 N$5945 N$5947 N$6024 N$6026 "Waveguide Crossing" sch_x=-102 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1584 N$5949 N$5951 N$6028 N$6030 "Waveguide Crossing" sch_x=-102 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1585 N$5953 N$5955 N$6032 N$6034 "Waveguide Crossing" sch_x=-102 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1586 N$5957 N$5959 N$6036 N$6821 "Waveguide Crossing" sch_x=-102 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1587 N$5961 N$5963 N$6745 N$6038 "Waveguide Crossing" sch_x=-100 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1588 N$5965 N$5967 N$6040 N$6042 "Waveguide Crossing" sch_x=-100 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1589 N$5969 N$5971 N$6044 N$6046 "Waveguide Crossing" sch_x=-100 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1590 N$5973 N$5975 N$6048 N$6050 "Waveguide Crossing" sch_x=-100 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1591 N$5977 N$5979 N$6052 N$6054 "Waveguide Crossing" sch_x=-100 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1592 N$5981 N$5983 N$6056 N$6058 "Waveguide Crossing" sch_x=-100 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1593 N$5985 N$5987 N$6060 N$6062 "Waveguide Crossing" sch_x=-100 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1594 N$5989 N$5991 N$6064 N$6066 "Waveguide Crossing" sch_x=-100 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1595 N$5993 N$5995 N$6068 N$6070 "Waveguide Crossing" sch_x=-100 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1596 N$5997 N$5999 N$6072 N$6074 "Waveguide Crossing" sch_x=-100 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1597 N$6001 N$6003 N$6076 N$6078 "Waveguide Crossing" sch_x=-100 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1598 N$6005 N$6007 N$6080 N$6082 "Waveguide Crossing" sch_x=-100 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1599 N$6009 N$6011 N$6084 N$6086 "Waveguide Crossing" sch_x=-100 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1600 N$6013 N$6015 N$6088 N$6090 "Waveguide Crossing" sch_x=-100 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1601 N$6017 N$6019 N$6092 N$6094 "Waveguide Crossing" sch_x=-100 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1602 N$6021 N$6023 N$6096 N$6098 "Waveguide Crossing" sch_x=-100 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1603 N$6025 N$6027 N$6100 N$6102 "Waveguide Crossing" sch_x=-100 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1604 N$6029 N$6031 N$6104 N$6106 "Waveguide Crossing" sch_x=-100 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1605 N$6033 N$6035 N$6108 N$6819 "Waveguide Crossing" sch_x=-100 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1606 N$6037 N$6039 N$6747 N$6110 "Waveguide Crossing" sch_x=-98 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1607 N$6041 N$6043 N$6112 N$6114 "Waveguide Crossing" sch_x=-98 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1608 N$6045 N$6047 N$6116 N$6118 "Waveguide Crossing" sch_x=-98 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1609 N$6049 N$6051 N$6120 N$6122 "Waveguide Crossing" sch_x=-98 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1610 N$6053 N$6055 N$6124 N$6126 "Waveguide Crossing" sch_x=-98 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1611 N$6057 N$6059 N$6128 N$6130 "Waveguide Crossing" sch_x=-98 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1612 N$6061 N$6063 N$6132 N$6134 "Waveguide Crossing" sch_x=-98 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1613 N$6065 N$6067 N$6136 N$6138 "Waveguide Crossing" sch_x=-98 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1614 N$6069 N$6071 N$6140 N$6142 "Waveguide Crossing" sch_x=-98 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1615 N$6073 N$6075 N$6144 N$6146 "Waveguide Crossing" sch_x=-98 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1616 N$6077 N$6079 N$6148 N$6150 "Waveguide Crossing" sch_x=-98 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1617 N$6081 N$6083 N$6152 N$6154 "Waveguide Crossing" sch_x=-98 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1618 N$6085 N$6087 N$6156 N$6158 "Waveguide Crossing" sch_x=-98 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1619 N$6089 N$6091 N$6160 N$6162 "Waveguide Crossing" sch_x=-98 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1620 N$6093 N$6095 N$6164 N$6166 "Waveguide Crossing" sch_x=-98 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1621 N$6097 N$6099 N$6168 N$6170 "Waveguide Crossing" sch_x=-98 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1622 N$6101 N$6103 N$6172 N$6174 "Waveguide Crossing" sch_x=-98 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1623 N$6105 N$6107 N$6176 N$6817 "Waveguide Crossing" sch_x=-98 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1624 N$6109 N$6111 N$6749 N$6178 "Waveguide Crossing" sch_x=-96 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1625 N$6113 N$6115 N$6180 N$6182 "Waveguide Crossing" sch_x=-96 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1626 N$6117 N$6119 N$6184 N$6186 "Waveguide Crossing" sch_x=-96 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1627 N$6121 N$6123 N$6188 N$6190 "Waveguide Crossing" sch_x=-96 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1628 N$6125 N$6127 N$6192 N$6194 "Waveguide Crossing" sch_x=-96 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1629 N$6129 N$6131 N$6196 N$6198 "Waveguide Crossing" sch_x=-96 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1630 N$6133 N$6135 N$6200 N$6202 "Waveguide Crossing" sch_x=-96 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1631 N$6137 N$6139 N$6204 N$6206 "Waveguide Crossing" sch_x=-96 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1632 N$6141 N$6143 N$6208 N$6210 "Waveguide Crossing" sch_x=-96 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1633 N$6145 N$6147 N$6212 N$6214 "Waveguide Crossing" sch_x=-96 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1634 N$6149 N$6151 N$6216 N$6218 "Waveguide Crossing" sch_x=-96 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1635 N$6153 N$6155 N$6220 N$6222 "Waveguide Crossing" sch_x=-96 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1636 N$6157 N$6159 N$6224 N$6226 "Waveguide Crossing" sch_x=-96 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1637 N$6161 N$6163 N$6228 N$6230 "Waveguide Crossing" sch_x=-96 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1638 N$6165 N$6167 N$6232 N$6234 "Waveguide Crossing" sch_x=-96 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1639 N$6169 N$6171 N$6236 N$6238 "Waveguide Crossing" sch_x=-96 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1640 N$6173 N$6175 N$6240 N$6815 "Waveguide Crossing" sch_x=-96 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1641 N$6177 N$6179 N$6751 N$6242 "Waveguide Crossing" sch_x=-94 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1642 N$6181 N$6183 N$6244 N$6246 "Waveguide Crossing" sch_x=-94 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1643 N$6185 N$6187 N$6248 N$6250 "Waveguide Crossing" sch_x=-94 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1644 N$6189 N$6191 N$6252 N$6254 "Waveguide Crossing" sch_x=-94 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1645 N$6193 N$6195 N$6256 N$6258 "Waveguide Crossing" sch_x=-94 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1646 N$6197 N$6199 N$6260 N$6262 "Waveguide Crossing" sch_x=-94 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1647 N$6201 N$6203 N$6264 N$6266 "Waveguide Crossing" sch_x=-94 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1648 N$6205 N$6207 N$6268 N$6270 "Waveguide Crossing" sch_x=-94 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1649 N$6209 N$6211 N$6272 N$6274 "Waveguide Crossing" sch_x=-94 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1650 N$6213 N$6215 N$6276 N$6278 "Waveguide Crossing" sch_x=-94 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1651 N$6217 N$6219 N$6280 N$6282 "Waveguide Crossing" sch_x=-94 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1652 N$6221 N$6223 N$6284 N$6286 "Waveguide Crossing" sch_x=-94 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1653 N$6225 N$6227 N$6288 N$6290 "Waveguide Crossing" sch_x=-94 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1654 N$6229 N$6231 N$6292 N$6294 "Waveguide Crossing" sch_x=-94 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1655 N$6233 N$6235 N$6296 N$6298 "Waveguide Crossing" sch_x=-94 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1656 N$6237 N$6239 N$6300 N$6813 "Waveguide Crossing" sch_x=-94 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1657 N$6241 N$6243 N$6753 N$6302 "Waveguide Crossing" sch_x=-92 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1658 N$6245 N$6247 N$6304 N$6306 "Waveguide Crossing" sch_x=-92 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1659 N$6249 N$6251 N$6308 N$6310 "Waveguide Crossing" sch_x=-92 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1660 N$6253 N$6255 N$6312 N$6314 "Waveguide Crossing" sch_x=-92 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1661 N$6257 N$6259 N$6316 N$6318 "Waveguide Crossing" sch_x=-92 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1662 N$6261 N$6263 N$6320 N$6322 "Waveguide Crossing" sch_x=-92 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1663 N$6265 N$6267 N$6324 N$6326 "Waveguide Crossing" sch_x=-92 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1664 N$6269 N$6271 N$6328 N$6330 "Waveguide Crossing" sch_x=-92 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1665 N$6273 N$6275 N$6332 N$6334 "Waveguide Crossing" sch_x=-92 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1666 N$6277 N$6279 N$6336 N$6338 "Waveguide Crossing" sch_x=-92 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1667 N$6281 N$6283 N$6340 N$6342 "Waveguide Crossing" sch_x=-92 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1668 N$6285 N$6287 N$6344 N$6346 "Waveguide Crossing" sch_x=-92 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1669 N$6289 N$6291 N$6348 N$6350 "Waveguide Crossing" sch_x=-92 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1670 N$6293 N$6295 N$6352 N$6354 "Waveguide Crossing" sch_x=-92 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1671 N$6297 N$6299 N$6356 N$6811 "Waveguide Crossing" sch_x=-92 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1672 N$6301 N$6303 N$6755 N$6358 "Waveguide Crossing" sch_x=-90 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1673 N$6305 N$6307 N$6360 N$6362 "Waveguide Crossing" sch_x=-90 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1674 N$6309 N$6311 N$6364 N$6366 "Waveguide Crossing" sch_x=-90 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1675 N$6313 N$6315 N$6368 N$6370 "Waveguide Crossing" sch_x=-90 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1676 N$6317 N$6319 N$6372 N$6374 "Waveguide Crossing" sch_x=-90 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1677 N$6321 N$6323 N$6376 N$6378 "Waveguide Crossing" sch_x=-90 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1678 N$6325 N$6327 N$6380 N$6382 "Waveguide Crossing" sch_x=-90 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1679 N$6329 N$6331 N$6384 N$6386 "Waveguide Crossing" sch_x=-90 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1680 N$6333 N$6335 N$6388 N$6390 "Waveguide Crossing" sch_x=-90 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1681 N$6337 N$6339 N$6392 N$6394 "Waveguide Crossing" sch_x=-90 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1682 N$6341 N$6343 N$6396 N$6398 "Waveguide Crossing" sch_x=-90 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1683 N$6345 N$6347 N$6400 N$6402 "Waveguide Crossing" sch_x=-90 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1684 N$6349 N$6351 N$6404 N$6406 "Waveguide Crossing" sch_x=-90 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1685 N$6353 N$6355 N$6408 N$6809 "Waveguide Crossing" sch_x=-90 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1686 N$6357 N$6359 N$6757 N$6410 "Waveguide Crossing" sch_x=-88 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1687 N$6361 N$6363 N$6412 N$6414 "Waveguide Crossing" sch_x=-88 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1688 N$6365 N$6367 N$6416 N$6418 "Waveguide Crossing" sch_x=-88 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1689 N$6369 N$6371 N$6420 N$6422 "Waveguide Crossing" sch_x=-88 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1690 N$6373 N$6375 N$6424 N$6426 "Waveguide Crossing" sch_x=-88 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1691 N$6377 N$6379 N$6428 N$6430 "Waveguide Crossing" sch_x=-88 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1692 N$6381 N$6383 N$6432 N$6434 "Waveguide Crossing" sch_x=-88 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1693 N$6385 N$6387 N$6436 N$6438 "Waveguide Crossing" sch_x=-88 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1694 N$6389 N$6391 N$6440 N$6442 "Waveguide Crossing" sch_x=-88 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1695 N$6393 N$6395 N$6444 N$6446 "Waveguide Crossing" sch_x=-88 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1696 N$6397 N$6399 N$6448 N$6450 "Waveguide Crossing" sch_x=-88 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1697 N$6401 N$6403 N$6452 N$6454 "Waveguide Crossing" sch_x=-88 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1698 N$6405 N$6407 N$6456 N$6807 "Waveguide Crossing" sch_x=-88 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1699 N$6409 N$6411 N$6759 N$6458 "Waveguide Crossing" sch_x=-86 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1700 N$6413 N$6415 N$6460 N$6462 "Waveguide Crossing" sch_x=-86 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1701 N$6417 N$6419 N$6464 N$6466 "Waveguide Crossing" sch_x=-86 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1702 N$6421 N$6423 N$6468 N$6470 "Waveguide Crossing" sch_x=-86 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1703 N$6425 N$6427 N$6472 N$6474 "Waveguide Crossing" sch_x=-86 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1704 N$6429 N$6431 N$6476 N$6478 "Waveguide Crossing" sch_x=-86 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1705 N$6433 N$6435 N$6480 N$6482 "Waveguide Crossing" sch_x=-86 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1706 N$6437 N$6439 N$6484 N$6486 "Waveguide Crossing" sch_x=-86 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1707 N$6441 N$6443 N$6488 N$6490 "Waveguide Crossing" sch_x=-86 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1708 N$6445 N$6447 N$6492 N$6494 "Waveguide Crossing" sch_x=-86 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1709 N$6449 N$6451 N$6496 N$6498 "Waveguide Crossing" sch_x=-86 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1710 N$6453 N$6455 N$6500 N$6805 "Waveguide Crossing" sch_x=-86 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1711 N$6457 N$6459 N$6761 N$6502 "Waveguide Crossing" sch_x=-84 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1712 N$6461 N$6463 N$6504 N$6506 "Waveguide Crossing" sch_x=-84 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1713 N$6465 N$6467 N$6508 N$6510 "Waveguide Crossing" sch_x=-84 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1714 N$6469 N$6471 N$6512 N$6514 "Waveguide Crossing" sch_x=-84 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1715 N$6473 N$6475 N$6516 N$6518 "Waveguide Crossing" sch_x=-84 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1716 N$6477 N$6479 N$6520 N$6522 "Waveguide Crossing" sch_x=-84 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1717 N$6481 N$6483 N$6524 N$6526 "Waveguide Crossing" sch_x=-84 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1718 N$6485 N$6487 N$6528 N$6530 "Waveguide Crossing" sch_x=-84 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1719 N$6489 N$6491 N$6532 N$6534 "Waveguide Crossing" sch_x=-84 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1720 N$6493 N$6495 N$6536 N$6538 "Waveguide Crossing" sch_x=-84 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1721 N$6497 N$6499 N$6540 N$6803 "Waveguide Crossing" sch_x=-84 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1722 N$6501 N$6503 N$6763 N$6542 "Waveguide Crossing" sch_x=-82 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1723 N$6505 N$6507 N$6544 N$6546 "Waveguide Crossing" sch_x=-82 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1724 N$6509 N$6511 N$6548 N$6550 "Waveguide Crossing" sch_x=-82 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1725 N$6513 N$6515 N$6552 N$6554 "Waveguide Crossing" sch_x=-82 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1726 N$6517 N$6519 N$6556 N$6558 "Waveguide Crossing" sch_x=-82 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1727 N$6521 N$6523 N$6560 N$6562 "Waveguide Crossing" sch_x=-82 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1728 N$6525 N$6527 N$6564 N$6566 "Waveguide Crossing" sch_x=-82 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1729 N$6529 N$6531 N$6568 N$6570 "Waveguide Crossing" sch_x=-82 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1730 N$6533 N$6535 N$6572 N$6574 "Waveguide Crossing" sch_x=-82 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1731 N$6537 N$6539 N$6576 N$6801 "Waveguide Crossing" sch_x=-82 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1732 N$6541 N$6543 N$6765 N$6578 "Waveguide Crossing" sch_x=-80 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1733 N$6545 N$6547 N$6580 N$6582 "Waveguide Crossing" sch_x=-80 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1734 N$6549 N$6551 N$6584 N$6586 "Waveguide Crossing" sch_x=-80 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1735 N$6553 N$6555 N$6588 N$6590 "Waveguide Crossing" sch_x=-80 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1736 N$6557 N$6559 N$6592 N$6594 "Waveguide Crossing" sch_x=-80 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1737 N$6561 N$6563 N$6596 N$6598 "Waveguide Crossing" sch_x=-80 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1738 N$6565 N$6567 N$6600 N$6602 "Waveguide Crossing" sch_x=-80 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1739 N$6569 N$6571 N$6604 N$6606 "Waveguide Crossing" sch_x=-80 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1740 N$6573 N$6575 N$6608 N$6799 "Waveguide Crossing" sch_x=-80 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1741 N$6577 N$6579 N$6767 N$6610 "Waveguide Crossing" sch_x=-78 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1742 N$6581 N$6583 N$6612 N$6614 "Waveguide Crossing" sch_x=-78 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1743 N$6585 N$6587 N$6616 N$6618 "Waveguide Crossing" sch_x=-78 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1744 N$6589 N$6591 N$6620 N$6622 "Waveguide Crossing" sch_x=-78 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1745 N$6593 N$6595 N$6624 N$6626 "Waveguide Crossing" sch_x=-78 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1746 N$6597 N$6599 N$6628 N$6630 "Waveguide Crossing" sch_x=-78 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1747 N$6601 N$6603 N$6632 N$6634 "Waveguide Crossing" sch_x=-78 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1748 N$6605 N$6607 N$6636 N$6797 "Waveguide Crossing" sch_x=-78 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1749 N$6609 N$6611 N$6769 N$6638 "Waveguide Crossing" sch_x=-76 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1750 N$6613 N$6615 N$6640 N$6642 "Waveguide Crossing" sch_x=-76 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1751 N$6617 N$6619 N$6644 N$6646 "Waveguide Crossing" sch_x=-76 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1752 N$6621 N$6623 N$6648 N$6650 "Waveguide Crossing" sch_x=-76 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1753 N$6625 N$6627 N$6652 N$6654 "Waveguide Crossing" sch_x=-76 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1754 N$6629 N$6631 N$6656 N$6658 "Waveguide Crossing" sch_x=-76 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1755 N$6633 N$6635 N$6660 N$6795 "Waveguide Crossing" sch_x=-76 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1756 N$6637 N$6639 N$6771 N$6662 "Waveguide Crossing" sch_x=-74 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1757 N$6641 N$6643 N$6664 N$6666 "Waveguide Crossing" sch_x=-74 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1758 N$6645 N$6647 N$6668 N$6670 "Waveguide Crossing" sch_x=-74 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1759 N$6649 N$6651 N$6672 N$6674 "Waveguide Crossing" sch_x=-74 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1760 N$6653 N$6655 N$6676 N$6678 "Waveguide Crossing" sch_x=-74 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1761 N$6657 N$6659 N$6680 N$6793 "Waveguide Crossing" sch_x=-74 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1762 N$6661 N$6663 N$6773 N$6682 "Waveguide Crossing" sch_x=-72 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1763 N$6665 N$6667 N$6684 N$6686 "Waveguide Crossing" sch_x=-72 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1764 N$6669 N$6671 N$6688 N$6690 "Waveguide Crossing" sch_x=-72 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1765 N$6673 N$6675 N$6692 N$6694 "Waveguide Crossing" sch_x=-72 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1766 N$6677 N$6679 N$6696 N$6791 "Waveguide Crossing" sch_x=-72 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1767 N$6681 N$6683 N$6775 N$6698 "Waveguide Crossing" sch_x=-70 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1768 N$6685 N$6687 N$6700 N$6702 "Waveguide Crossing" sch_x=-70 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1769 N$6689 N$6691 N$6704 N$6706 "Waveguide Crossing" sch_x=-70 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1770 N$6693 N$6695 N$6708 N$6789 "Waveguide Crossing" sch_x=-70 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1771 N$6697 N$6699 N$6777 N$6710 "Waveguide Crossing" sch_x=-68 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1772 N$6701 N$6703 N$6712 N$6714 "Waveguide Crossing" sch_x=-68 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1773 N$6705 N$6707 N$6716 N$6787 "Waveguide Crossing" sch_x=-68 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1774 N$6709 N$6711 N$6779 N$6718 "Waveguide Crossing" sch_x=-66 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1775 N$6713 N$6715 N$6720 N$6785 "Waveguide Crossing" sch_x=-66 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1776 N$6717 N$6719 N$6781 N$6783 "Waveguide Crossing" sch_x=-64 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S977 N$6784 N$6786 N$4189 N$3650 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S978 N$6788 N$6790 N$3652 N$3654 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S979 N$6792 N$6794 N$3656 N$3658 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S980 N$6796 N$6798 N$3660 N$3662 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S981 N$6800 N$6802 N$3664 N$3666 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S982 N$6804 N$6806 N$3668 N$3670 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S983 N$6808 N$6810 N$3672 N$3674 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S984 N$6812 N$6814 N$3676 N$3678 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S985 N$6816 N$6818 N$3680 N$3682 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S986 N$6820 N$6822 N$3684 N$3686 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S987 N$6824 N$6826 N$3688 N$3690 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S988 N$6828 N$6830 N$3692 N$3694 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S989 N$6832 N$6834 N$3696 N$3698 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S990 N$6836 N$6838 N$3700 N$3702 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S991 N$6840 N$6842 N$3704 N$3706 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S992 N$6844 N$6848 N$3708 N$4191 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C993 N$3649 N$3651 N$4129 N$3710 "Waveguide Crossing" sch_x=-60 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C994 N$3653 N$3655 N$3712 N$3714 "Waveguide Crossing" sch_x=-60 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C995 N$3657 N$3659 N$3716 N$3718 "Waveguide Crossing" sch_x=-60 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C996 N$3661 N$3663 N$3720 N$3722 "Waveguide Crossing" sch_x=-60 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C997 N$3665 N$3667 N$3724 N$3726 "Waveguide Crossing" sch_x=-60 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C998 N$3669 N$3671 N$3728 N$3730 "Waveguide Crossing" sch_x=-60 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C999 N$3673 N$3675 N$3732 N$3734 "Waveguide Crossing" sch_x=-60 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1000 N$3677 N$3679 N$3736 N$3738 "Waveguide Crossing" sch_x=-60 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1001 N$3681 N$3683 N$3740 N$3742 "Waveguide Crossing" sch_x=-60 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1002 N$3685 N$3687 N$3744 N$3746 "Waveguide Crossing" sch_x=-60 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1003 N$3689 N$3691 N$3748 N$3750 "Waveguide Crossing" sch_x=-60 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1004 N$3693 N$3695 N$3752 N$3754 "Waveguide Crossing" sch_x=-60 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1005 N$3697 N$3699 N$3756 N$3758 "Waveguide Crossing" sch_x=-60 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1006 N$3701 N$3703 N$3760 N$3762 "Waveguide Crossing" sch_x=-60 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1007 N$3705 N$3707 N$3764 N$4187 "Waveguide Crossing" sch_x=-60 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1008 N$3709 N$3711 N$4131 N$3766 "Waveguide Crossing" sch_x=-58 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1009 N$3713 N$3715 N$3768 N$3770 "Waveguide Crossing" sch_x=-58 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1010 N$3717 N$3719 N$3772 N$3774 "Waveguide Crossing" sch_x=-58 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1011 N$3721 N$3723 N$3776 N$3778 "Waveguide Crossing" sch_x=-58 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1012 N$3725 N$3727 N$3780 N$3782 "Waveguide Crossing" sch_x=-58 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1013 N$3729 N$3731 N$3784 N$3786 "Waveguide Crossing" sch_x=-58 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1014 N$3733 N$3735 N$3788 N$3790 "Waveguide Crossing" sch_x=-58 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1015 N$3737 N$3739 N$3792 N$3794 "Waveguide Crossing" sch_x=-58 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1016 N$3741 N$3743 N$3796 N$3798 "Waveguide Crossing" sch_x=-58 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1017 N$3745 N$3747 N$3800 N$3802 "Waveguide Crossing" sch_x=-58 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1018 N$3749 N$3751 N$3804 N$3806 "Waveguide Crossing" sch_x=-58 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1019 N$3753 N$3755 N$3808 N$3810 "Waveguide Crossing" sch_x=-58 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1020 N$3757 N$3759 N$3812 N$3814 "Waveguide Crossing" sch_x=-58 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1021 N$3761 N$3763 N$3816 N$4185 "Waveguide Crossing" sch_x=-58 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1022 N$3765 N$3767 N$4133 N$3818 "Waveguide Crossing" sch_x=-56 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1023 N$3769 N$3771 N$3820 N$3822 "Waveguide Crossing" sch_x=-56 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1024 N$3773 N$3775 N$3824 N$3826 "Waveguide Crossing" sch_x=-56 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1025 N$3777 N$3779 N$3828 N$3830 "Waveguide Crossing" sch_x=-56 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1026 N$3781 N$3783 N$3832 N$3834 "Waveguide Crossing" sch_x=-56 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1027 N$3785 N$3787 N$3836 N$3838 "Waveguide Crossing" sch_x=-56 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1028 N$3789 N$3791 N$3840 N$3842 "Waveguide Crossing" sch_x=-56 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1029 N$3793 N$3795 N$3844 N$3846 "Waveguide Crossing" sch_x=-56 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1030 N$3797 N$3799 N$3848 N$3850 "Waveguide Crossing" sch_x=-56 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1031 N$3801 N$3803 N$3852 N$3854 "Waveguide Crossing" sch_x=-56 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1032 N$3805 N$3807 N$3856 N$3858 "Waveguide Crossing" sch_x=-56 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1033 N$3809 N$3811 N$3860 N$3862 "Waveguide Crossing" sch_x=-56 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1034 N$3813 N$3815 N$3864 N$4183 "Waveguide Crossing" sch_x=-56 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1035 N$3817 N$3819 N$4135 N$3866 "Waveguide Crossing" sch_x=-54 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1036 N$3821 N$3823 N$3868 N$3870 "Waveguide Crossing" sch_x=-54 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1037 N$3825 N$3827 N$3872 N$3874 "Waveguide Crossing" sch_x=-54 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1038 N$3829 N$3831 N$3876 N$3878 "Waveguide Crossing" sch_x=-54 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1039 N$3833 N$3835 N$3880 N$3882 "Waveguide Crossing" sch_x=-54 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1040 N$3837 N$3839 N$3884 N$3886 "Waveguide Crossing" sch_x=-54 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1041 N$3841 N$3843 N$3888 N$3890 "Waveguide Crossing" sch_x=-54 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1042 N$3845 N$3847 N$3892 N$3894 "Waveguide Crossing" sch_x=-54 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1043 N$3849 N$3851 N$3896 N$3898 "Waveguide Crossing" sch_x=-54 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1044 N$3853 N$3855 N$3900 N$3902 "Waveguide Crossing" sch_x=-54 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1045 N$3857 N$3859 N$3904 N$3906 "Waveguide Crossing" sch_x=-54 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1046 N$3861 N$3863 N$3908 N$4181 "Waveguide Crossing" sch_x=-54 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1047 N$3865 N$3867 N$4137 N$3910 "Waveguide Crossing" sch_x=-52 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1048 N$3869 N$3871 N$3912 N$3914 "Waveguide Crossing" sch_x=-52 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1049 N$3873 N$3875 N$3916 N$3918 "Waveguide Crossing" sch_x=-52 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1050 N$3877 N$3879 N$3920 N$3922 "Waveguide Crossing" sch_x=-52 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1051 N$3881 N$3883 N$3924 N$3926 "Waveguide Crossing" sch_x=-52 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1052 N$3885 N$3887 N$3928 N$3930 "Waveguide Crossing" sch_x=-52 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1053 N$3889 N$3891 N$3932 N$3934 "Waveguide Crossing" sch_x=-52 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1054 N$3893 N$3895 N$3936 N$3938 "Waveguide Crossing" sch_x=-52 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1055 N$3897 N$3899 N$3940 N$3942 "Waveguide Crossing" sch_x=-52 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1056 N$3901 N$3903 N$3944 N$3946 "Waveguide Crossing" sch_x=-52 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1057 N$3905 N$3907 N$3948 N$4179 "Waveguide Crossing" sch_x=-52 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1058 N$3909 N$3911 N$4139 N$3950 "Waveguide Crossing" sch_x=-50 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1059 N$3913 N$3915 N$3952 N$3954 "Waveguide Crossing" sch_x=-50 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1060 N$3917 N$3919 N$3956 N$3958 "Waveguide Crossing" sch_x=-50 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1061 N$3921 N$3923 N$3960 N$3962 "Waveguide Crossing" sch_x=-50 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1062 N$3925 N$3927 N$3964 N$3966 "Waveguide Crossing" sch_x=-50 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1063 N$3929 N$3931 N$3968 N$3970 "Waveguide Crossing" sch_x=-50 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1064 N$3933 N$3935 N$3972 N$3974 "Waveguide Crossing" sch_x=-50 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1065 N$3937 N$3939 N$3976 N$3978 "Waveguide Crossing" sch_x=-50 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1066 N$3941 N$3943 N$3980 N$3982 "Waveguide Crossing" sch_x=-50 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1067 N$3945 N$3947 N$3984 N$4177 "Waveguide Crossing" sch_x=-50 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1068 N$3949 N$3951 N$4141 N$3986 "Waveguide Crossing" sch_x=-48 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1069 N$3953 N$3955 N$3988 N$3990 "Waveguide Crossing" sch_x=-48 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1070 N$3957 N$3959 N$3992 N$3994 "Waveguide Crossing" sch_x=-48 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1071 N$3961 N$3963 N$3996 N$3998 "Waveguide Crossing" sch_x=-48 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1072 N$3965 N$3967 N$4000 N$4002 "Waveguide Crossing" sch_x=-48 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1073 N$3969 N$3971 N$4004 N$4006 "Waveguide Crossing" sch_x=-48 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1074 N$3973 N$3975 N$4008 N$4010 "Waveguide Crossing" sch_x=-48 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1075 N$3977 N$3979 N$4012 N$4014 "Waveguide Crossing" sch_x=-48 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1076 N$3981 N$3983 N$4016 N$4175 "Waveguide Crossing" sch_x=-48 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1077 N$3985 N$3987 N$4143 N$4018 "Waveguide Crossing" sch_x=-46 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1078 N$3989 N$3991 N$4020 N$4022 "Waveguide Crossing" sch_x=-46 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1079 N$3993 N$3995 N$4024 N$4026 "Waveguide Crossing" sch_x=-46 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1080 N$3997 N$3999 N$4028 N$4030 "Waveguide Crossing" sch_x=-46 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1081 N$4001 N$4003 N$4032 N$4034 "Waveguide Crossing" sch_x=-46 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1082 N$4005 N$4007 N$4036 N$4038 "Waveguide Crossing" sch_x=-46 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1083 N$4009 N$4011 N$4040 N$4042 "Waveguide Crossing" sch_x=-46 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1084 N$4013 N$4015 N$4044 N$4173 "Waveguide Crossing" sch_x=-46 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1085 N$4017 N$4019 N$4145 N$4046 "Waveguide Crossing" sch_x=-44 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1086 N$4021 N$4023 N$4048 N$4050 "Waveguide Crossing" sch_x=-44 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1087 N$4025 N$4027 N$4052 N$4054 "Waveguide Crossing" sch_x=-44 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1088 N$4029 N$4031 N$4056 N$4058 "Waveguide Crossing" sch_x=-44 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1089 N$4033 N$4035 N$4060 N$4062 "Waveguide Crossing" sch_x=-44 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1090 N$4037 N$4039 N$4064 N$4066 "Waveguide Crossing" sch_x=-44 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1091 N$4041 N$4043 N$4068 N$4171 "Waveguide Crossing" sch_x=-44 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1092 N$4045 N$4047 N$4147 N$4070 "Waveguide Crossing" sch_x=-42 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1093 N$4049 N$4051 N$4072 N$4074 "Waveguide Crossing" sch_x=-42 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1094 N$4053 N$4055 N$4076 N$4078 "Waveguide Crossing" sch_x=-42 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1095 N$4057 N$4059 N$4080 N$4082 "Waveguide Crossing" sch_x=-42 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1096 N$4061 N$4063 N$4084 N$4086 "Waveguide Crossing" sch_x=-42 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1097 N$4065 N$4067 N$4088 N$4169 "Waveguide Crossing" sch_x=-42 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1098 N$4069 N$4071 N$4149 N$4090 "Waveguide Crossing" sch_x=-40 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1099 N$4073 N$4075 N$4092 N$4094 "Waveguide Crossing" sch_x=-40 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1100 N$4077 N$4079 N$4096 N$4098 "Waveguide Crossing" sch_x=-40 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1101 N$4081 N$4083 N$4100 N$4102 "Waveguide Crossing" sch_x=-40 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1102 N$4085 N$4087 N$4104 N$4167 "Waveguide Crossing" sch_x=-40 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1103 N$4089 N$4091 N$4151 N$4106 "Waveguide Crossing" sch_x=-38 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1104 N$4093 N$4095 N$4108 N$4110 "Waveguide Crossing" sch_x=-38 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1105 N$4097 N$4099 N$4112 N$4114 "Waveguide Crossing" sch_x=-38 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1106 N$4101 N$4103 N$4116 N$4165 "Waveguide Crossing" sch_x=-38 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1107 N$4105 N$4107 N$4153 N$4118 "Waveguide Crossing" sch_x=-36 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1108 N$4109 N$4111 N$4120 N$4122 "Waveguide Crossing" sch_x=-36 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1109 N$4113 N$4115 N$4124 N$4163 "Waveguide Crossing" sch_x=-36 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1110 N$4117 N$4119 N$4155 N$4126 "Waveguide Crossing" sch_x=-34 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1111 N$4121 N$4123 N$4128 N$4161 "Waveguide Crossing" sch_x=-34 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1112 N$4125 N$4127 N$4157 N$4159 "Waveguide Crossing" sch_x=-32 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S905 N$4160 N$4162 N$3501 N$3362 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S906 N$4164 N$4166 N$3364 N$3366 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S907 N$4168 N$4170 N$3368 N$3370 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S908 N$4172 N$4174 N$3372 N$3374 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S909 N$4176 N$4178 N$3376 N$3378 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S910 N$4180 N$4182 N$3380 N$3382 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S911 N$4184 N$4186 N$3384 N$3386 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S912 N$4188 N$4192 N$3388 N$3503 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C913 N$3361 N$3363 N$3473 N$3390 "Waveguide Crossing" sch_x=-28 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C914 N$3365 N$3367 N$3392 N$3394 "Waveguide Crossing" sch_x=-28 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C915 N$3369 N$3371 N$3396 N$3398 "Waveguide Crossing" sch_x=-28 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C916 N$3373 N$3375 N$3400 N$3402 "Waveguide Crossing" sch_x=-28 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C917 N$3377 N$3379 N$3404 N$3406 "Waveguide Crossing" sch_x=-28 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C918 N$3381 N$3383 N$3408 N$3410 "Waveguide Crossing" sch_x=-28 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C919 N$3385 N$3387 N$3412 N$3499 "Waveguide Crossing" sch_x=-28 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C920 N$3389 N$3391 N$3475 N$3414 "Waveguide Crossing" sch_x=-26 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C921 N$3393 N$3395 N$3416 N$3418 "Waveguide Crossing" sch_x=-26 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C922 N$3397 N$3399 N$3420 N$3422 "Waveguide Crossing" sch_x=-26 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C923 N$3401 N$3403 N$3424 N$3426 "Waveguide Crossing" sch_x=-26 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C924 N$3405 N$3407 N$3428 N$3430 "Waveguide Crossing" sch_x=-26 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C925 N$3409 N$3411 N$3432 N$3497 "Waveguide Crossing" sch_x=-26 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C926 N$3413 N$3415 N$3477 N$3434 "Waveguide Crossing" sch_x=-24 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C927 N$3417 N$3419 N$3436 N$3438 "Waveguide Crossing" sch_x=-24 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C928 N$3421 N$3423 N$3440 N$3442 "Waveguide Crossing" sch_x=-24 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C929 N$3425 N$3427 N$3444 N$3446 "Waveguide Crossing" sch_x=-24 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C930 N$3429 N$3431 N$3448 N$3495 "Waveguide Crossing" sch_x=-24 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C931 N$3433 N$3435 N$3479 N$3450 "Waveguide Crossing" sch_x=-22 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C932 N$3437 N$3439 N$3452 N$3454 "Waveguide Crossing" sch_x=-22 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C933 N$3441 N$3443 N$3456 N$3458 "Waveguide Crossing" sch_x=-22 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C934 N$3445 N$3447 N$3460 N$3493 "Waveguide Crossing" sch_x=-22 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C935 N$3449 N$3451 N$3481 N$3462 "Waveguide Crossing" sch_x=-20 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C936 N$3453 N$3455 N$3464 N$3466 "Waveguide Crossing" sch_x=-20 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C937 N$3457 N$3459 N$3468 N$3491 "Waveguide Crossing" sch_x=-20 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C938 N$3461 N$3463 N$3483 N$3470 "Waveguide Crossing" sch_x=-18 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C939 N$3465 N$3467 N$3472 N$3489 "Waveguide Crossing" sch_x=-18 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C940 N$3469 N$3471 N$3485 N$3487 "Waveguide Crossing" sch_x=-16 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S885 N$3488 N$3490 N$3317 N$3282 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S886 N$3492 N$3494 N$3284 N$3286 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S887 N$3496 N$3498 N$3288 N$3290 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S888 N$3500 N$3504 N$3292 N$3319 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C889 N$3281 N$3283 N$3305 N$3294 "Waveguide Crossing" sch_x=-12 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C890 N$3285 N$3287 N$3296 N$3298 "Waveguide Crossing" sch_x=-12 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C891 N$3289 N$3291 N$3300 N$3315 "Waveguide Crossing" sch_x=-12 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C892 N$3293 N$3295 N$3307 N$3302 "Waveguide Crossing" sch_x=-10 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C893 N$3297 N$3299 N$3304 N$3313 "Waveguide Crossing" sch_x=-10 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C894 N$3301 N$3303 N$3309 N$3311 "Waveguide Crossing" sch_x=-8 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S833 N$3502 N$3474 N$3141 N$3106 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S834 N$3476 N$3478 N$3108 N$3110 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S835 N$3480 N$3482 N$3112 N$3114 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S836 N$3484 N$3486 N$3116 N$3143 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C837 N$3105 N$3107 N$3129 N$3118 "Waveguide Crossing" sch_x=-12 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C838 N$3109 N$3111 N$3120 N$3122 "Waveguide Crossing" sch_x=-12 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C839 N$3113 N$3115 N$3124 N$3139 "Waveguide Crossing" sch_x=-12 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C840 N$3117 N$3119 N$3131 N$3126 "Waveguide Crossing" sch_x=-10 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C841 N$3121 N$3123 N$3128 N$3137 "Waveguide Crossing" sch_x=-10 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C842 N$3125 N$3127 N$3133 N$3135 "Waveguide Crossing" sch_x=-8 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S729 N$4190 N$4130 N$2861 N$2722 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S730 N$4132 N$4134 N$2724 N$2726 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S731 N$4136 N$4138 N$2728 N$2730 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S732 N$4140 N$4142 N$2732 N$2734 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S733 N$4144 N$4146 N$2736 N$2738 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S734 N$4148 N$4150 N$2740 N$2742 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S735 N$4152 N$4154 N$2744 N$2746 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S736 N$4156 N$4158 N$2748 N$2863 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C737 N$2721 N$2723 N$2833 N$2750 "Waveguide Crossing" sch_x=-28 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C738 N$2725 N$2727 N$2752 N$2754 "Waveguide Crossing" sch_x=-28 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C739 N$2729 N$2731 N$2756 N$2758 "Waveguide Crossing" sch_x=-28 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C740 N$2733 N$2735 N$2760 N$2762 "Waveguide Crossing" sch_x=-28 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C741 N$2737 N$2739 N$2764 N$2766 "Waveguide Crossing" sch_x=-28 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C742 N$2741 N$2743 N$2768 N$2770 "Waveguide Crossing" sch_x=-28 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C743 N$2745 N$2747 N$2772 N$2859 "Waveguide Crossing" sch_x=-28 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C744 N$2749 N$2751 N$2835 N$2774 "Waveguide Crossing" sch_x=-26 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C745 N$2753 N$2755 N$2776 N$2778 "Waveguide Crossing" sch_x=-26 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C746 N$2757 N$2759 N$2780 N$2782 "Waveguide Crossing" sch_x=-26 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C747 N$2761 N$2763 N$2784 N$2786 "Waveguide Crossing" sch_x=-26 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C748 N$2765 N$2767 N$2788 N$2790 "Waveguide Crossing" sch_x=-26 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C749 N$2769 N$2771 N$2792 N$2857 "Waveguide Crossing" sch_x=-26 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C750 N$2773 N$2775 N$2837 N$2794 "Waveguide Crossing" sch_x=-24 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C751 N$2777 N$2779 N$2796 N$2798 "Waveguide Crossing" sch_x=-24 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C752 N$2781 N$2783 N$2800 N$2802 "Waveguide Crossing" sch_x=-24 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C753 N$2785 N$2787 N$2804 N$2806 "Waveguide Crossing" sch_x=-24 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C754 N$2789 N$2791 N$2808 N$2855 "Waveguide Crossing" sch_x=-24 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C755 N$2793 N$2795 N$2839 N$2810 "Waveguide Crossing" sch_x=-22 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C756 N$2797 N$2799 N$2812 N$2814 "Waveguide Crossing" sch_x=-22 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C757 N$2801 N$2803 N$2816 N$2818 "Waveguide Crossing" sch_x=-22 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C758 N$2805 N$2807 N$2820 N$2853 "Waveguide Crossing" sch_x=-22 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C759 N$2809 N$2811 N$2841 N$2822 "Waveguide Crossing" sch_x=-20 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C760 N$2813 N$2815 N$2824 N$2826 "Waveguide Crossing" sch_x=-20 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C761 N$2817 N$2819 N$2828 N$2851 "Waveguide Crossing" sch_x=-20 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C762 N$2821 N$2823 N$2843 N$2830 "Waveguide Crossing" sch_x=-18 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C763 N$2825 N$2827 N$2832 N$2849 "Waveguide Crossing" sch_x=-18 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C764 N$2829 N$2831 N$2845 N$2847 "Waveguide Crossing" sch_x=-16 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S709 N$2848 N$2850 N$2677 N$2642 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S710 N$2852 N$2854 N$2644 N$2646 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S711 N$2856 N$2858 N$2648 N$2650 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S712 N$2860 N$2864 N$2652 N$2679 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C713 N$2641 N$2643 N$2665 N$2654 "Waveguide Crossing" sch_x=-12 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C714 N$2645 N$2647 N$2656 N$2658 "Waveguide Crossing" sch_x=-12 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C715 N$2649 N$2651 N$2660 N$2675 "Waveguide Crossing" sch_x=-12 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C716 N$2653 N$2655 N$2667 N$2662 "Waveguide Crossing" sch_x=-10 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C717 N$2657 N$2659 N$2664 N$2673 "Waveguide Crossing" sch_x=-10 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C718 N$2661 N$2663 N$2669 N$2671 "Waveguide Crossing" sch_x=-8 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S657 N$2862 N$2834 N$2501 N$2466 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S658 N$2836 N$2838 N$2468 N$2470 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S659 N$2840 N$2842 N$2472 N$2474 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S660 N$2844 N$2846 N$2476 N$2503 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C661 N$2465 N$2467 N$2489 N$2478 "Waveguide Crossing" sch_x=-12 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C662 N$2469 N$2471 N$2480 N$2482 "Waveguide Crossing" sch_x=-12 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C663 N$2473 N$2475 N$2484 N$2499 "Waveguide Crossing" sch_x=-12 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C664 N$2477 N$2479 N$2491 N$2486 "Waveguide Crossing" sch_x=-10 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C665 N$2481 N$2483 N$2488 N$2497 "Waveguide Crossing" sch_x=-10 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C666 N$2485 N$2487 N$2493 N$2495 "Waveguide Crossing" sch_x=-8 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S353 N$6846 N$6722 N$1821 N$1282 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S354 N$6724 N$6726 N$1284 N$1286 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S355 N$6728 N$6730 N$1288 N$1290 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S356 N$6732 N$6734 N$1292 N$1294 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S357 N$6736 N$6738 N$1296 N$1298 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S358 N$6740 N$6742 N$1300 N$1302 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S359 N$6744 N$6746 N$1304 N$1306 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S360 N$6748 N$6750 N$1308 N$1310 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S361 N$6752 N$6754 N$1312 N$1314 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S362 N$6756 N$6758 N$1316 N$1318 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S363 N$6760 N$6762 N$1320 N$1322 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S364 N$6764 N$6766 N$1324 N$1326 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S365 N$6768 N$6770 N$1328 N$1330 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S366 N$6772 N$6774 N$1332 N$1334 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S367 N$6776 N$6778 N$1336 N$1338 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S368 N$6780 N$6782 N$1340 N$1823 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C369 N$1281 N$1283 N$1761 N$1342 "Waveguide Crossing" sch_x=-60 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C370 N$1285 N$1287 N$1344 N$1346 "Waveguide Crossing" sch_x=-60 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C371 N$1289 N$1291 N$1348 N$1350 "Waveguide Crossing" sch_x=-60 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C372 N$1293 N$1295 N$1352 N$1354 "Waveguide Crossing" sch_x=-60 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C373 N$1297 N$1299 N$1356 N$1358 "Waveguide Crossing" sch_x=-60 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C374 N$1301 N$1303 N$1360 N$1362 "Waveguide Crossing" sch_x=-60 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C375 N$1305 N$1307 N$1364 N$1366 "Waveguide Crossing" sch_x=-60 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C376 N$1309 N$1311 N$1368 N$1370 "Waveguide Crossing" sch_x=-60 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C377 N$1313 N$1315 N$1372 N$1374 "Waveguide Crossing" sch_x=-60 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C378 N$1317 N$1319 N$1376 N$1378 "Waveguide Crossing" sch_x=-60 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C379 N$1321 N$1323 N$1380 N$1382 "Waveguide Crossing" sch_x=-60 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C380 N$1325 N$1327 N$1384 N$1386 "Waveguide Crossing" sch_x=-60 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C381 N$1329 N$1331 N$1388 N$1390 "Waveguide Crossing" sch_x=-60 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C382 N$1333 N$1335 N$1392 N$1394 "Waveguide Crossing" sch_x=-60 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C383 N$1337 N$1339 N$1396 N$1819 "Waveguide Crossing" sch_x=-60 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C384 N$1341 N$1343 N$1763 N$1398 "Waveguide Crossing" sch_x=-58 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C385 N$1345 N$1347 N$1400 N$1402 "Waveguide Crossing" sch_x=-58 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C386 N$1349 N$1351 N$1404 N$1406 "Waveguide Crossing" sch_x=-58 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C387 N$1353 N$1355 N$1408 N$1410 "Waveguide Crossing" sch_x=-58 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C388 N$1357 N$1359 N$1412 N$1414 "Waveguide Crossing" sch_x=-58 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C389 N$1361 N$1363 N$1416 N$1418 "Waveguide Crossing" sch_x=-58 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C390 N$1365 N$1367 N$1420 N$1422 "Waveguide Crossing" sch_x=-58 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C391 N$1369 N$1371 N$1424 N$1426 "Waveguide Crossing" sch_x=-58 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C392 N$1373 N$1375 N$1428 N$1430 "Waveguide Crossing" sch_x=-58 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C393 N$1377 N$1379 N$1432 N$1434 "Waveguide Crossing" sch_x=-58 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C394 N$1381 N$1383 N$1436 N$1438 "Waveguide Crossing" sch_x=-58 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C395 N$1385 N$1387 N$1440 N$1442 "Waveguide Crossing" sch_x=-58 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C396 N$1389 N$1391 N$1444 N$1446 "Waveguide Crossing" sch_x=-58 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C397 N$1393 N$1395 N$1448 N$1817 "Waveguide Crossing" sch_x=-58 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C398 N$1397 N$1399 N$1765 N$1450 "Waveguide Crossing" sch_x=-56 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C399 N$1401 N$1403 N$1452 N$1454 "Waveguide Crossing" sch_x=-56 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C400 N$1405 N$1407 N$1456 N$1458 "Waveguide Crossing" sch_x=-56 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C401 N$1409 N$1411 N$1460 N$1462 "Waveguide Crossing" sch_x=-56 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C402 N$1413 N$1415 N$1464 N$1466 "Waveguide Crossing" sch_x=-56 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C403 N$1417 N$1419 N$1468 N$1470 "Waveguide Crossing" sch_x=-56 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C404 N$1421 N$1423 N$1472 N$1474 "Waveguide Crossing" sch_x=-56 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C405 N$1425 N$1427 N$1476 N$1478 "Waveguide Crossing" sch_x=-56 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C406 N$1429 N$1431 N$1480 N$1482 "Waveguide Crossing" sch_x=-56 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C407 N$1433 N$1435 N$1484 N$1486 "Waveguide Crossing" sch_x=-56 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C408 N$1437 N$1439 N$1488 N$1490 "Waveguide Crossing" sch_x=-56 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C409 N$1441 N$1443 N$1492 N$1494 "Waveguide Crossing" sch_x=-56 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C410 N$1445 N$1447 N$1496 N$1815 "Waveguide Crossing" sch_x=-56 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C411 N$1449 N$1451 N$1767 N$1498 "Waveguide Crossing" sch_x=-54 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C412 N$1453 N$1455 N$1500 N$1502 "Waveguide Crossing" sch_x=-54 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C413 N$1457 N$1459 N$1504 N$1506 "Waveguide Crossing" sch_x=-54 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C414 N$1461 N$1463 N$1508 N$1510 "Waveguide Crossing" sch_x=-54 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C415 N$1465 N$1467 N$1512 N$1514 "Waveguide Crossing" sch_x=-54 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C416 N$1469 N$1471 N$1516 N$1518 "Waveguide Crossing" sch_x=-54 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C417 N$1473 N$1475 N$1520 N$1522 "Waveguide Crossing" sch_x=-54 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C418 N$1477 N$1479 N$1524 N$1526 "Waveguide Crossing" sch_x=-54 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C419 N$1481 N$1483 N$1528 N$1530 "Waveguide Crossing" sch_x=-54 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C420 N$1485 N$1487 N$1532 N$1534 "Waveguide Crossing" sch_x=-54 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C421 N$1489 N$1491 N$1536 N$1538 "Waveguide Crossing" sch_x=-54 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C422 N$1493 N$1495 N$1540 N$1813 "Waveguide Crossing" sch_x=-54 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C423 N$1497 N$1499 N$1769 N$1542 "Waveguide Crossing" sch_x=-52 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C424 N$1501 N$1503 N$1544 N$1546 "Waveguide Crossing" sch_x=-52 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C425 N$1505 N$1507 N$1548 N$1550 "Waveguide Crossing" sch_x=-52 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C426 N$1509 N$1511 N$1552 N$1554 "Waveguide Crossing" sch_x=-52 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C427 N$1513 N$1515 N$1556 N$1558 "Waveguide Crossing" sch_x=-52 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C428 N$1517 N$1519 N$1560 N$1562 "Waveguide Crossing" sch_x=-52 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C429 N$1521 N$1523 N$1564 N$1566 "Waveguide Crossing" sch_x=-52 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C430 N$1525 N$1527 N$1568 N$1570 "Waveguide Crossing" sch_x=-52 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C431 N$1529 N$1531 N$1572 N$1574 "Waveguide Crossing" sch_x=-52 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C432 N$1533 N$1535 N$1576 N$1578 "Waveguide Crossing" sch_x=-52 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C433 N$1537 N$1539 N$1580 N$1811 "Waveguide Crossing" sch_x=-52 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C434 N$1541 N$1543 N$1771 N$1582 "Waveguide Crossing" sch_x=-50 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C435 N$1545 N$1547 N$1584 N$1586 "Waveguide Crossing" sch_x=-50 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C436 N$1549 N$1551 N$1588 N$1590 "Waveguide Crossing" sch_x=-50 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C437 N$1553 N$1555 N$1592 N$1594 "Waveguide Crossing" sch_x=-50 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C438 N$1557 N$1559 N$1596 N$1598 "Waveguide Crossing" sch_x=-50 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C439 N$1561 N$1563 N$1600 N$1602 "Waveguide Crossing" sch_x=-50 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C440 N$1565 N$1567 N$1604 N$1606 "Waveguide Crossing" sch_x=-50 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C441 N$1569 N$1571 N$1608 N$1610 "Waveguide Crossing" sch_x=-50 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C442 N$1573 N$1575 N$1612 N$1614 "Waveguide Crossing" sch_x=-50 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C443 N$1577 N$1579 N$1616 N$1809 "Waveguide Crossing" sch_x=-50 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C444 N$1581 N$1583 N$1773 N$1618 "Waveguide Crossing" sch_x=-48 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C445 N$1585 N$1587 N$1620 N$1622 "Waveguide Crossing" sch_x=-48 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C446 N$1589 N$1591 N$1624 N$1626 "Waveguide Crossing" sch_x=-48 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C447 N$1593 N$1595 N$1628 N$1630 "Waveguide Crossing" sch_x=-48 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C448 N$1597 N$1599 N$1632 N$1634 "Waveguide Crossing" sch_x=-48 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C449 N$1601 N$1603 N$1636 N$1638 "Waveguide Crossing" sch_x=-48 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C450 N$1605 N$1607 N$1640 N$1642 "Waveguide Crossing" sch_x=-48 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C451 N$1609 N$1611 N$1644 N$1646 "Waveguide Crossing" sch_x=-48 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C452 N$1613 N$1615 N$1648 N$1807 "Waveguide Crossing" sch_x=-48 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C453 N$1617 N$1619 N$1775 N$1650 "Waveguide Crossing" sch_x=-46 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C454 N$1621 N$1623 N$1652 N$1654 "Waveguide Crossing" sch_x=-46 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C455 N$1625 N$1627 N$1656 N$1658 "Waveguide Crossing" sch_x=-46 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C456 N$1629 N$1631 N$1660 N$1662 "Waveguide Crossing" sch_x=-46 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C457 N$1633 N$1635 N$1664 N$1666 "Waveguide Crossing" sch_x=-46 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C458 N$1637 N$1639 N$1668 N$1670 "Waveguide Crossing" sch_x=-46 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C459 N$1641 N$1643 N$1672 N$1674 "Waveguide Crossing" sch_x=-46 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C460 N$1645 N$1647 N$1676 N$1805 "Waveguide Crossing" sch_x=-46 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C461 N$1649 N$1651 N$1777 N$1678 "Waveguide Crossing" sch_x=-44 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C462 N$1653 N$1655 N$1680 N$1682 "Waveguide Crossing" sch_x=-44 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C463 N$1657 N$1659 N$1684 N$1686 "Waveguide Crossing" sch_x=-44 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C464 N$1661 N$1663 N$1688 N$1690 "Waveguide Crossing" sch_x=-44 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C465 N$1665 N$1667 N$1692 N$1694 "Waveguide Crossing" sch_x=-44 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C466 N$1669 N$1671 N$1696 N$1698 "Waveguide Crossing" sch_x=-44 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C467 N$1673 N$1675 N$1700 N$1803 "Waveguide Crossing" sch_x=-44 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C468 N$1677 N$1679 N$1779 N$1702 "Waveguide Crossing" sch_x=-42 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C469 N$1681 N$1683 N$1704 N$1706 "Waveguide Crossing" sch_x=-42 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C470 N$1685 N$1687 N$1708 N$1710 "Waveguide Crossing" sch_x=-42 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C471 N$1689 N$1691 N$1712 N$1714 "Waveguide Crossing" sch_x=-42 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C472 N$1693 N$1695 N$1716 N$1718 "Waveguide Crossing" sch_x=-42 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C473 N$1697 N$1699 N$1720 N$1801 "Waveguide Crossing" sch_x=-42 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C474 N$1701 N$1703 N$1781 N$1722 "Waveguide Crossing" sch_x=-40 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C475 N$1705 N$1707 N$1724 N$1726 "Waveguide Crossing" sch_x=-40 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C476 N$1709 N$1711 N$1728 N$1730 "Waveguide Crossing" sch_x=-40 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C477 N$1713 N$1715 N$1732 N$1734 "Waveguide Crossing" sch_x=-40 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C478 N$1717 N$1719 N$1736 N$1799 "Waveguide Crossing" sch_x=-40 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C479 N$1721 N$1723 N$1783 N$1738 "Waveguide Crossing" sch_x=-38 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C480 N$1725 N$1727 N$1740 N$1742 "Waveguide Crossing" sch_x=-38 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C481 N$1729 N$1731 N$1744 N$1746 "Waveguide Crossing" sch_x=-38 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C482 N$1733 N$1735 N$1748 N$1797 "Waveguide Crossing" sch_x=-38 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C483 N$1737 N$1739 N$1785 N$1750 "Waveguide Crossing" sch_x=-36 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C484 N$1741 N$1743 N$1752 N$1754 "Waveguide Crossing" sch_x=-36 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C485 N$1745 N$1747 N$1756 N$1795 "Waveguide Crossing" sch_x=-36 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C486 N$1749 N$1751 N$1787 N$1758 "Waveguide Crossing" sch_x=-34 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C487 N$1753 N$1755 N$1760 N$1793 "Waveguide Crossing" sch_x=-34 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C488 N$1757 N$1759 N$1789 N$1791 "Waveguide Crossing" sch_x=-32 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S281 N$1792 N$1794 N$1133 N$994 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S282 N$1796 N$1798 N$996 N$998 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S283 N$1800 N$1802 N$1000 N$1002 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S284 N$1804 N$1806 N$1004 N$1006 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S285 N$1808 N$1810 N$1008 N$1010 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S286 N$1812 N$1814 N$1012 N$1014 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S287 N$1816 N$1818 N$1016 N$1018 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S288 N$1820 N$1824 N$1020 N$1135 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C289 N$993 N$995 N$1105 N$1022 "Waveguide Crossing" sch_x=-28 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C290 N$997 N$999 N$1024 N$1026 "Waveguide Crossing" sch_x=-28 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C291 N$1001 N$1003 N$1028 N$1030 "Waveguide Crossing" sch_x=-28 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C292 N$1005 N$1007 N$1032 N$1034 "Waveguide Crossing" sch_x=-28 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C293 N$1009 N$1011 N$1036 N$1038 "Waveguide Crossing" sch_x=-28 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C294 N$1013 N$1015 N$1040 N$1042 "Waveguide Crossing" sch_x=-28 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C295 N$1017 N$1019 N$1044 N$1131 "Waveguide Crossing" sch_x=-28 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C296 N$1021 N$1023 N$1107 N$1046 "Waveguide Crossing" sch_x=-26 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C297 N$1025 N$1027 N$1048 N$1050 "Waveguide Crossing" sch_x=-26 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C298 N$1029 N$1031 N$1052 N$1054 "Waveguide Crossing" sch_x=-26 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C299 N$1033 N$1035 N$1056 N$1058 "Waveguide Crossing" sch_x=-26 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C300 N$1037 N$1039 N$1060 N$1062 "Waveguide Crossing" sch_x=-26 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C301 N$1041 N$1043 N$1064 N$1129 "Waveguide Crossing" sch_x=-26 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C302 N$1045 N$1047 N$1109 N$1066 "Waveguide Crossing" sch_x=-24 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C303 N$1049 N$1051 N$1068 N$1070 "Waveguide Crossing" sch_x=-24 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C304 N$1053 N$1055 N$1072 N$1074 "Waveguide Crossing" sch_x=-24 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C305 N$1057 N$1059 N$1076 N$1078 "Waveguide Crossing" sch_x=-24 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C306 N$1061 N$1063 N$1080 N$1127 "Waveguide Crossing" sch_x=-24 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C307 N$1065 N$1067 N$1111 N$1082 "Waveguide Crossing" sch_x=-22 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C308 N$1069 N$1071 N$1084 N$1086 "Waveguide Crossing" sch_x=-22 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C309 N$1073 N$1075 N$1088 N$1090 "Waveguide Crossing" sch_x=-22 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C310 N$1077 N$1079 N$1092 N$1125 "Waveguide Crossing" sch_x=-22 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C311 N$1081 N$1083 N$1113 N$1094 "Waveguide Crossing" sch_x=-20 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C312 N$1085 N$1087 N$1096 N$1098 "Waveguide Crossing" sch_x=-20 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C313 N$1089 N$1091 N$1100 N$1123 "Waveguide Crossing" sch_x=-20 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C314 N$1093 N$1095 N$1115 N$1102 "Waveguide Crossing" sch_x=-18 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C315 N$1097 N$1099 N$1104 N$1121 "Waveguide Crossing" sch_x=-18 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C316 N$1101 N$1103 N$1117 N$1119 "Waveguide Crossing" sch_x=-16 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S261 N$1120 N$1122 N$949 N$914 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S262 N$1124 N$1126 N$916 N$918 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S263 N$1128 N$1130 N$920 N$922 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S264 N$1132 N$1136 N$924 N$951 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C265 N$913 N$915 N$937 N$926 "Waveguide Crossing" sch_x=-12 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C266 N$917 N$919 N$928 N$930 "Waveguide Crossing" sch_x=-12 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C267 N$921 N$923 N$932 N$947 "Waveguide Crossing" sch_x=-12 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C268 N$925 N$927 N$939 N$934 "Waveguide Crossing" sch_x=-10 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C269 N$929 N$931 N$936 N$945 "Waveguide Crossing" sch_x=-10 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C270 N$933 N$935 N$941 N$943 "Waveguide Crossing" sch_x=-8 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S209 N$1134 N$1106 N$773 N$738 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S210 N$1108 N$1110 N$740 N$742 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S211 N$1112 N$1114 N$744 N$746 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S212 N$1116 N$1118 N$748 N$775 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C213 N$737 N$739 N$761 N$750 "Waveguide Crossing" sch_x=-12 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C214 N$741 N$743 N$752 N$754 "Waveguide Crossing" sch_x=-12 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C215 N$745 N$747 N$756 N$771 "Waveguide Crossing" sch_x=-12 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C216 N$749 N$751 N$763 N$758 "Waveguide Crossing" sch_x=-10 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C217 N$753 N$755 N$760 N$769 "Waveguide Crossing" sch_x=-10 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C218 N$757 N$759 N$765 N$767 "Waveguide Crossing" sch_x=-8 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S105 N$1822 N$1762 N$493 N$354 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S106 N$1764 N$1766 N$356 N$358 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S107 N$1768 N$1770 N$360 N$362 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S108 N$1772 N$1774 N$364 N$366 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S109 N$1776 N$1778 N$368 N$370 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S110 N$1780 N$1782 N$372 N$374 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S111 N$1784 N$1786 N$376 N$378 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S112 N$1788 N$1790 N$380 N$495 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C113 N$353 N$355 N$465 N$382 "Waveguide Crossing" sch_x=-28 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C114 N$357 N$359 N$384 N$386 "Waveguide Crossing" sch_x=-28 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C115 N$361 N$363 N$388 N$390 "Waveguide Crossing" sch_x=-28 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C116 N$365 N$367 N$392 N$394 "Waveguide Crossing" sch_x=-28 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C117 N$369 N$371 N$396 N$398 "Waveguide Crossing" sch_x=-28 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C118 N$373 N$375 N$400 N$402 "Waveguide Crossing" sch_x=-28 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C119 N$377 N$379 N$404 N$491 "Waveguide Crossing" sch_x=-28 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C120 N$381 N$383 N$467 N$406 "Waveguide Crossing" sch_x=-26 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C121 N$385 N$387 N$408 N$410 "Waveguide Crossing" sch_x=-26 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C122 N$389 N$391 N$412 N$414 "Waveguide Crossing" sch_x=-26 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C123 N$393 N$395 N$416 N$418 "Waveguide Crossing" sch_x=-26 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C124 N$397 N$399 N$420 N$422 "Waveguide Crossing" sch_x=-26 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C125 N$401 N$403 N$424 N$489 "Waveguide Crossing" sch_x=-26 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C126 N$405 N$407 N$469 N$426 "Waveguide Crossing" sch_x=-24 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C127 N$409 N$411 N$428 N$430 "Waveguide Crossing" sch_x=-24 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C128 N$413 N$415 N$432 N$434 "Waveguide Crossing" sch_x=-24 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C129 N$417 N$419 N$436 N$438 "Waveguide Crossing" sch_x=-24 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C130 N$421 N$423 N$440 N$487 "Waveguide Crossing" sch_x=-24 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C131 N$425 N$427 N$471 N$442 "Waveguide Crossing" sch_x=-22 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C132 N$429 N$431 N$444 N$446 "Waveguide Crossing" sch_x=-22 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C133 N$433 N$435 N$448 N$450 "Waveguide Crossing" sch_x=-22 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C134 N$437 N$439 N$452 N$485 "Waveguide Crossing" sch_x=-22 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C135 N$441 N$443 N$473 N$454 "Waveguide Crossing" sch_x=-20 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C136 N$445 N$447 N$456 N$458 "Waveguide Crossing" sch_x=-20 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C137 N$449 N$451 N$460 N$483 "Waveguide Crossing" sch_x=-20 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C138 N$453 N$455 N$475 N$462 "Waveguide Crossing" sch_x=-18 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C139 N$457 N$459 N$464 N$481 "Waveguide Crossing" sch_x=-18 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C140 N$461 N$463 N$477 N$479 "Waveguide Crossing" sch_x=-16 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S85 N$480 N$482 N$309 N$274 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S86 N$484 N$486 N$276 N$278 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S87 N$488 N$490 N$280 N$282 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S88 N$492 N$496 N$284 N$311 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C89 N$273 N$275 N$297 N$286 "Waveguide Crossing" sch_x=-12 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C90 N$277 N$279 N$288 N$290 "Waveguide Crossing" sch_x=-12 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C91 N$281 N$283 N$292 N$307 "Waveguide Crossing" sch_x=-12 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C92 N$285 N$287 N$299 N$294 "Waveguide Crossing" sch_x=-10 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C93 N$289 N$291 N$296 N$305 "Waveguide Crossing" sch_x=-10 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C94 N$293 N$295 N$301 N$303 "Waveguide Crossing" sch_x=-8 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S33 N$494 N$466 N$133 N$98 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S34 N$468 N$470 N$100 N$102 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S35 N$472 N$474 N$104 N$106 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S36 N$476 N$478 N$108 N$135 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C37 N$97 N$99 N$121 N$110 "Waveguide Crossing" sch_x=-12 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C38 N$101 N$103 N$112 N$114 "Waveguide Crossing" sch_x=-12 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C39 N$105 N$107 N$116 N$131 "Waveguide Crossing" sch_x=-12 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C40 N$109 N$111 N$123 N$118 "Waveguide Crossing" sch_x=-10 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C41 N$113 N$115 N$120 N$129 "Waveguide Crossing" sch_x=-10 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C42 N$117 N$119 N$125 N$127 "Waveguide Crossing" sch_x=-8 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1 N$134 N$122 N$1 N$3 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=62.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2 N$124 N$126 N$5 N$11 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=61.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3 N$34689 N$2 N$13 N$15 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=63.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4 N$8 N$34690 N$17 N$23 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S5 N$34691 N$10 N$25 N$27 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6 N$12 N$34692 N$29 N$35 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S7 N$14 N$22 N$37 N$34693 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=63.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S8 N$20 N$24 N$34694 N$39 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S9 N$26 N$34 N$41 N$34695 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S10 N$32 N$36 N$34696 N$47 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S11 N$38 N$46 N$174 N$162 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=62.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S12 N$44 N$48 N$164 N$166 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=61.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C13 N$4 N$6 N$7 N$9 "Waveguide Crossing" sch_x=-4 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C14 N$16 N$18 N$21 N$19 "Waveguide Crossing" sch_x=0 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C15 N$28 N$30 N$33 N$31 "Waveguide Crossing" sch_x=0 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C16 N$40 N$42 N$45 N$43 "Waveguide Crossing" sch_x=4 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S17 N$128 N$130 N$49 N$51 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=58.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S18 N$132 N$136 N$53 N$59 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=57.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S19 N$34697 N$50 N$61 N$63 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S20 N$56 N$34698 N$65 N$71 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S21 N$34699 N$58 N$73 N$75 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S22 N$60 N$34700 N$77 N$83 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S23 N$62 N$70 N$85 N$34701 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S24 N$68 N$72 N$34702 N$87 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S25 N$74 N$82 N$89 N$34703 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S26 N$80 N$84 N$34704 N$95 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S27 N$86 N$94 N$168 N$170 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=58.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S28 N$92 N$96 N$172 N$176 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=57.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C29 N$52 N$54 N$55 N$57 "Waveguide Crossing" sch_x=-4 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C30 N$64 N$66 N$69 N$67 "Waveguide Crossing" sch_x=0 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C31 N$76 N$78 N$81 N$79 "Waveguide Crossing" sch_x=0 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C32 N$88 N$90 N$93 N$91 "Waveguide Crossing" sch_x=4 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C47 N$161 N$150 N$137 N$139 "Waveguide Crossing" sch_x=12 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C48 N$152 N$154 N$141 N$143 "Waveguide Crossing" sch_x=12 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C49 N$156 N$171 N$145 N$147 "Waveguide Crossing" sch_x=12 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C50 N$163 N$158 N$149 N$151 "Waveguide Crossing" sch_x=10 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C51 N$160 N$169 N$153 N$155 "Waveguide Crossing" sch_x=10 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C52 N$165 N$167 N$157 N$159 "Waveguide Crossing" sch_x=8 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S43 N$173 N$138 N$638 N$610 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S44 N$140 N$142 N$612 N$614 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S45 N$144 N$146 N$616 N$618 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S46 N$148 N$175 N$620 N$622 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S53 N$310 N$298 N$177 N$179 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=54.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S54 N$300 N$302 N$181 N$187 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=53.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S55 N$34705 N$178 N$189 N$191 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S56 N$184 N$34706 N$193 N$199 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S57 N$34707 N$186 N$201 N$203 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S58 N$188 N$34708 N$205 N$211 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S59 N$190 N$198 N$213 N$34709 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S60 N$196 N$200 N$34710 N$215 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S61 N$202 N$210 N$217 N$34711 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S62 N$208 N$212 N$34712 N$223 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S63 N$214 N$222 N$350 N$338 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=54.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S64 N$220 N$224 N$340 N$342 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=53.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C65 N$180 N$182 N$183 N$185 "Waveguide Crossing" sch_x=-4 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C66 N$192 N$194 N$197 N$195 "Waveguide Crossing" sch_x=0 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C67 N$204 N$206 N$209 N$207 "Waveguide Crossing" sch_x=0 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C68 N$216 N$218 N$221 N$219 "Waveguide Crossing" sch_x=4 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S69 N$304 N$306 N$225 N$227 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=50.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S70 N$308 N$312 N$229 N$235 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=49.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S71 N$34713 N$226 N$237 N$239 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S72 N$232 N$34714 N$241 N$247 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S73 N$34715 N$234 N$249 N$251 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S74 N$236 N$34716 N$253 N$259 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S75 N$238 N$246 N$261 N$34717 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S76 N$244 N$248 N$34718 N$263 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S77 N$250 N$258 N$265 N$34719 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S78 N$256 N$260 N$34720 N$271 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S79 N$262 N$270 N$344 N$346 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=50.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S80 N$268 N$272 N$348 N$352 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=49.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C81 N$228 N$230 N$231 N$233 "Waveguide Crossing" sch_x=-4 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C82 N$240 N$242 N$245 N$243 "Waveguide Crossing" sch_x=0 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C83 N$252 N$254 N$257 N$255 "Waveguide Crossing" sch_x=0 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C84 N$264 N$266 N$269 N$267 "Waveguide Crossing" sch_x=4 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C99 N$337 N$326 N$313 N$315 "Waveguide Crossing" sch_x=12 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C100 N$328 N$330 N$317 N$319 "Waveguide Crossing" sch_x=12 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C101 N$332 N$347 N$321 N$323 "Waveguide Crossing" sch_x=12 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C102 N$339 N$334 N$325 N$327 "Waveguide Crossing" sch_x=10 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C103 N$336 N$345 N$329 N$331 "Waveguide Crossing" sch_x=10 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C104 N$341 N$343 N$333 N$335 "Waveguide Crossing" sch_x=8 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S95 N$349 N$314 N$624 N$626 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S96 N$316 N$318 N$628 N$630 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S97 N$320 N$322 N$632 N$634 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S98 N$324 N$351 N$636 N$640 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C149 N$609 N$526 N$497 N$499 "Waveguide Crossing" sch_x=28 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C150 N$528 N$530 N$501 N$503 "Waveguide Crossing" sch_x=28 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C151 N$532 N$534 N$505 N$507 "Waveguide Crossing" sch_x=28 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C152 N$536 N$538 N$509 N$511 "Waveguide Crossing" sch_x=28 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C153 N$540 N$542 N$513 N$515 "Waveguide Crossing" sch_x=28 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C154 N$544 N$546 N$517 N$519 "Waveguide Crossing" sch_x=28 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C155 N$548 N$635 N$521 N$523 "Waveguide Crossing" sch_x=28 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C156 N$611 N$550 N$525 N$527 "Waveguide Crossing" sch_x=26 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C157 N$552 N$554 N$529 N$531 "Waveguide Crossing" sch_x=26 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C158 N$556 N$558 N$533 N$535 "Waveguide Crossing" sch_x=26 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C159 N$560 N$562 N$537 N$539 "Waveguide Crossing" sch_x=26 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C160 N$564 N$566 N$541 N$543 "Waveguide Crossing" sch_x=26 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C161 N$568 N$633 N$545 N$547 "Waveguide Crossing" sch_x=26 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C162 N$613 N$570 N$549 N$551 "Waveguide Crossing" sch_x=24 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C163 N$572 N$574 N$553 N$555 "Waveguide Crossing" sch_x=24 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C164 N$576 N$578 N$557 N$559 "Waveguide Crossing" sch_x=24 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C165 N$580 N$582 N$561 N$563 "Waveguide Crossing" sch_x=24 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C166 N$584 N$631 N$565 N$567 "Waveguide Crossing" sch_x=24 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C167 N$615 N$586 N$569 N$571 "Waveguide Crossing" sch_x=22 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C168 N$588 N$590 N$573 N$575 "Waveguide Crossing" sch_x=22 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C169 N$592 N$594 N$577 N$579 "Waveguide Crossing" sch_x=22 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C170 N$596 N$629 N$581 N$583 "Waveguide Crossing" sch_x=22 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C171 N$617 N$598 N$585 N$587 "Waveguide Crossing" sch_x=20 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C172 N$600 N$602 N$589 N$591 "Waveguide Crossing" sch_x=20 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C173 N$604 N$627 N$593 N$595 "Waveguide Crossing" sch_x=20 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C174 N$619 N$606 N$597 N$599 "Waveguide Crossing" sch_x=18 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C175 N$608 N$625 N$601 N$603 "Waveguide Crossing" sch_x=18 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C176 N$621 N$623 N$605 N$607 "Waveguide Crossing" sch_x=16 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S141 N$637 N$498 N$2366 N$2306 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S142 N$500 N$502 N$2308 N$2310 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S143 N$504 N$506 N$2312 N$2314 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S144 N$508 N$510 N$2316 N$2318 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S145 N$512 N$514 N$2320 N$2322 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S146 N$516 N$518 N$2324 N$2326 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S147 N$520 N$522 N$2328 N$2330 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S148 N$524 N$639 N$2332 N$2334 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S177 N$774 N$762 N$641 N$643 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=46.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S178 N$764 N$766 N$645 N$651 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=45.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S179 N$34721 N$642 N$653 N$655 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S180 N$648 N$34722 N$657 N$663 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S181 N$34723 N$650 N$665 N$667 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S182 N$652 N$34724 N$669 N$675 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S183 N$654 N$662 N$677 N$34725 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S184 N$660 N$664 N$34726 N$679 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S185 N$666 N$674 N$681 N$34727 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S186 N$672 N$676 N$34728 N$687 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S187 N$678 N$686 N$814 N$802 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=46.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S188 N$684 N$688 N$804 N$806 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=45.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C189 N$644 N$646 N$647 N$649 "Waveguide Crossing" sch_x=-4 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C190 N$656 N$658 N$661 N$659 "Waveguide Crossing" sch_x=0 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C191 N$668 N$670 N$673 N$671 "Waveguide Crossing" sch_x=0 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C192 N$680 N$682 N$685 N$683 "Waveguide Crossing" sch_x=4 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S193 N$768 N$770 N$689 N$691 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=42.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S194 N$772 N$776 N$693 N$699 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=41.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S195 N$34729 N$690 N$701 N$703 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S196 N$696 N$34730 N$705 N$711 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S197 N$34731 N$698 N$713 N$715 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S198 N$700 N$34732 N$717 N$723 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S199 N$702 N$710 N$725 N$34733 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S200 N$708 N$712 N$34734 N$727 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S201 N$714 N$722 N$729 N$34735 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S202 N$720 N$724 N$34736 N$735 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S203 N$726 N$734 N$808 N$810 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=42.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S204 N$732 N$736 N$812 N$816 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=41.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C205 N$692 N$694 N$695 N$697 "Waveguide Crossing" sch_x=-4 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C206 N$704 N$706 N$709 N$707 "Waveguide Crossing" sch_x=0 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C207 N$716 N$718 N$721 N$719 "Waveguide Crossing" sch_x=0 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C208 N$728 N$730 N$733 N$731 "Waveguide Crossing" sch_x=4 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C223 N$801 N$790 N$777 N$779 "Waveguide Crossing" sch_x=12 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C224 N$792 N$794 N$781 N$783 "Waveguide Crossing" sch_x=12 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C225 N$796 N$811 N$785 N$787 "Waveguide Crossing" sch_x=12 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C226 N$803 N$798 N$789 N$791 "Waveguide Crossing" sch_x=10 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C227 N$800 N$809 N$793 N$795 "Waveguide Crossing" sch_x=10 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C228 N$805 N$807 N$797 N$799 "Waveguide Crossing" sch_x=8 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S219 N$813 N$778 N$1278 N$1250 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S220 N$780 N$782 N$1252 N$1254 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S221 N$784 N$786 N$1256 N$1258 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S222 N$788 N$815 N$1260 N$1262 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S229 N$950 N$938 N$817 N$819 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=38.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S230 N$940 N$942 N$821 N$827 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=37.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S231 N$34737 N$818 N$829 N$831 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S232 N$824 N$34738 N$833 N$839 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S233 N$34739 N$826 N$841 N$843 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S234 N$828 N$34740 N$845 N$851 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S235 N$830 N$838 N$853 N$34741 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S236 N$836 N$840 N$34742 N$855 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S237 N$842 N$850 N$857 N$34743 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S238 N$848 N$852 N$34744 N$863 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S239 N$854 N$862 N$990 N$978 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=38.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S240 N$860 N$864 N$980 N$982 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=37.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C241 N$820 N$822 N$823 N$825 "Waveguide Crossing" sch_x=-4 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C242 N$832 N$834 N$837 N$835 "Waveguide Crossing" sch_x=0 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C243 N$844 N$846 N$849 N$847 "Waveguide Crossing" sch_x=0 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C244 N$856 N$858 N$861 N$859 "Waveguide Crossing" sch_x=4 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S245 N$944 N$946 N$865 N$867 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=34.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S246 N$948 N$952 N$869 N$875 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=33.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S247 N$34745 N$866 N$877 N$879 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S248 N$872 N$34746 N$881 N$887 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S249 N$34747 N$874 N$889 N$891 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S250 N$876 N$34748 N$893 N$899 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S251 N$878 N$886 N$901 N$34749 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S252 N$884 N$888 N$34750 N$903 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S253 N$890 N$898 N$905 N$34751 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S254 N$896 N$900 N$34752 N$911 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S255 N$902 N$910 N$984 N$986 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=34.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S256 N$908 N$912 N$988 N$992 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=33.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C257 N$868 N$870 N$871 N$873 "Waveguide Crossing" sch_x=-4 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C258 N$880 N$882 N$885 N$883 "Waveguide Crossing" sch_x=0 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C259 N$892 N$894 N$897 N$895 "Waveguide Crossing" sch_x=0 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C260 N$904 N$906 N$909 N$907 "Waveguide Crossing" sch_x=4 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C275 N$977 N$966 N$953 N$955 "Waveguide Crossing" sch_x=12 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C276 N$968 N$970 N$957 N$959 "Waveguide Crossing" sch_x=12 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C277 N$972 N$987 N$961 N$963 "Waveguide Crossing" sch_x=12 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C278 N$979 N$974 N$965 N$967 "Waveguide Crossing" sch_x=10 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C279 N$976 N$985 N$969 N$971 "Waveguide Crossing" sch_x=10 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C280 N$981 N$983 N$973 N$975 "Waveguide Crossing" sch_x=8 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S271 N$989 N$954 N$1264 N$1266 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S272 N$956 N$958 N$1268 N$1270 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S273 N$960 N$962 N$1272 N$1274 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S274 N$964 N$991 N$1276 N$1280 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C325 N$1249 N$1166 N$1137 N$1139 "Waveguide Crossing" sch_x=28 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C326 N$1168 N$1170 N$1141 N$1143 "Waveguide Crossing" sch_x=28 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C327 N$1172 N$1174 N$1145 N$1147 "Waveguide Crossing" sch_x=28 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C328 N$1176 N$1178 N$1149 N$1151 "Waveguide Crossing" sch_x=28 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C329 N$1180 N$1182 N$1153 N$1155 "Waveguide Crossing" sch_x=28 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C330 N$1184 N$1186 N$1157 N$1159 "Waveguide Crossing" sch_x=28 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C331 N$1188 N$1275 N$1161 N$1163 "Waveguide Crossing" sch_x=28 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C332 N$1251 N$1190 N$1165 N$1167 "Waveguide Crossing" sch_x=26 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C333 N$1192 N$1194 N$1169 N$1171 "Waveguide Crossing" sch_x=26 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C334 N$1196 N$1198 N$1173 N$1175 "Waveguide Crossing" sch_x=26 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C335 N$1200 N$1202 N$1177 N$1179 "Waveguide Crossing" sch_x=26 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C336 N$1204 N$1206 N$1181 N$1183 "Waveguide Crossing" sch_x=26 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C337 N$1208 N$1273 N$1185 N$1187 "Waveguide Crossing" sch_x=26 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C338 N$1253 N$1210 N$1189 N$1191 "Waveguide Crossing" sch_x=24 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C339 N$1212 N$1214 N$1193 N$1195 "Waveguide Crossing" sch_x=24 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C340 N$1216 N$1218 N$1197 N$1199 "Waveguide Crossing" sch_x=24 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C341 N$1220 N$1222 N$1201 N$1203 "Waveguide Crossing" sch_x=24 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C342 N$1224 N$1271 N$1205 N$1207 "Waveguide Crossing" sch_x=24 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C343 N$1255 N$1226 N$1209 N$1211 "Waveguide Crossing" sch_x=22 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C344 N$1228 N$1230 N$1213 N$1215 "Waveguide Crossing" sch_x=22 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C345 N$1232 N$1234 N$1217 N$1219 "Waveguide Crossing" sch_x=22 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C346 N$1236 N$1269 N$1221 N$1223 "Waveguide Crossing" sch_x=22 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C347 N$1257 N$1238 N$1225 N$1227 "Waveguide Crossing" sch_x=20 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C348 N$1240 N$1242 N$1229 N$1231 "Waveguide Crossing" sch_x=20 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C349 N$1244 N$1267 N$1233 N$1235 "Waveguide Crossing" sch_x=20 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C350 N$1259 N$1246 N$1237 N$1239 "Waveguide Crossing" sch_x=18 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C351 N$1248 N$1265 N$1241 N$1243 "Waveguide Crossing" sch_x=18 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C352 N$1261 N$1263 N$1245 N$1247 "Waveguide Crossing" sch_x=16 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S317 N$1277 N$1138 N$2336 N$2338 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S318 N$1140 N$1142 N$2340 N$2342 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S319 N$1144 N$1146 N$2344 N$2346 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S320 N$1148 N$1150 N$2348 N$2350 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S321 N$1152 N$1154 N$2352 N$2354 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S322 N$1156 N$1158 N$2356 N$2358 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S323 N$1160 N$1162 N$2360 N$2362 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S324 N$1164 N$1279 N$2364 N$2368 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C505 N$2305 N$1886 N$1825 N$1827 "Waveguide Crossing" sch_x=60 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C506 N$1888 N$1890 N$1829 N$1831 "Waveguide Crossing" sch_x=60 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C507 N$1892 N$1894 N$1833 N$1835 "Waveguide Crossing" sch_x=60 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C508 N$1896 N$1898 N$1837 N$1839 "Waveguide Crossing" sch_x=60 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C509 N$1900 N$1902 N$1841 N$1843 "Waveguide Crossing" sch_x=60 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C510 N$1904 N$1906 N$1845 N$1847 "Waveguide Crossing" sch_x=60 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C511 N$1908 N$1910 N$1849 N$1851 "Waveguide Crossing" sch_x=60 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C512 N$1912 N$1914 N$1853 N$1855 "Waveguide Crossing" sch_x=60 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C513 N$1916 N$1918 N$1857 N$1859 "Waveguide Crossing" sch_x=60 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C514 N$1920 N$1922 N$1861 N$1863 "Waveguide Crossing" sch_x=60 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C515 N$1924 N$1926 N$1865 N$1867 "Waveguide Crossing" sch_x=60 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C516 N$1928 N$1930 N$1869 N$1871 "Waveguide Crossing" sch_x=60 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C517 N$1932 N$1934 N$1873 N$1875 "Waveguide Crossing" sch_x=60 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C518 N$1936 N$1938 N$1877 N$1879 "Waveguide Crossing" sch_x=60 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C519 N$1940 N$2363 N$1881 N$1883 "Waveguide Crossing" sch_x=60 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C520 N$2307 N$1942 N$1885 N$1887 "Waveguide Crossing" sch_x=58 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C521 N$1944 N$1946 N$1889 N$1891 "Waveguide Crossing" sch_x=58 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C522 N$1948 N$1950 N$1893 N$1895 "Waveguide Crossing" sch_x=58 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C523 N$1952 N$1954 N$1897 N$1899 "Waveguide Crossing" sch_x=58 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C524 N$1956 N$1958 N$1901 N$1903 "Waveguide Crossing" sch_x=58 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C525 N$1960 N$1962 N$1905 N$1907 "Waveguide Crossing" sch_x=58 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C526 N$1964 N$1966 N$1909 N$1911 "Waveguide Crossing" sch_x=58 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C527 N$1968 N$1970 N$1913 N$1915 "Waveguide Crossing" sch_x=58 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C528 N$1972 N$1974 N$1917 N$1919 "Waveguide Crossing" sch_x=58 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C529 N$1976 N$1978 N$1921 N$1923 "Waveguide Crossing" sch_x=58 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C530 N$1980 N$1982 N$1925 N$1927 "Waveguide Crossing" sch_x=58 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C531 N$1984 N$1986 N$1929 N$1931 "Waveguide Crossing" sch_x=58 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C532 N$1988 N$1990 N$1933 N$1935 "Waveguide Crossing" sch_x=58 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C533 N$1992 N$2361 N$1937 N$1939 "Waveguide Crossing" sch_x=58 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C534 N$2309 N$1994 N$1941 N$1943 "Waveguide Crossing" sch_x=56 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C535 N$1996 N$1998 N$1945 N$1947 "Waveguide Crossing" sch_x=56 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C536 N$2000 N$2002 N$1949 N$1951 "Waveguide Crossing" sch_x=56 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C537 N$2004 N$2006 N$1953 N$1955 "Waveguide Crossing" sch_x=56 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C538 N$2008 N$2010 N$1957 N$1959 "Waveguide Crossing" sch_x=56 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C539 N$2012 N$2014 N$1961 N$1963 "Waveguide Crossing" sch_x=56 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C540 N$2016 N$2018 N$1965 N$1967 "Waveguide Crossing" sch_x=56 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C541 N$2020 N$2022 N$1969 N$1971 "Waveguide Crossing" sch_x=56 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C542 N$2024 N$2026 N$1973 N$1975 "Waveguide Crossing" sch_x=56 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C543 N$2028 N$2030 N$1977 N$1979 "Waveguide Crossing" sch_x=56 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C544 N$2032 N$2034 N$1981 N$1983 "Waveguide Crossing" sch_x=56 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C545 N$2036 N$2038 N$1985 N$1987 "Waveguide Crossing" sch_x=56 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C546 N$2040 N$2359 N$1989 N$1991 "Waveguide Crossing" sch_x=56 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C547 N$2311 N$2042 N$1993 N$1995 "Waveguide Crossing" sch_x=54 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C548 N$2044 N$2046 N$1997 N$1999 "Waveguide Crossing" sch_x=54 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C549 N$2048 N$2050 N$2001 N$2003 "Waveguide Crossing" sch_x=54 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C550 N$2052 N$2054 N$2005 N$2007 "Waveguide Crossing" sch_x=54 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C551 N$2056 N$2058 N$2009 N$2011 "Waveguide Crossing" sch_x=54 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C552 N$2060 N$2062 N$2013 N$2015 "Waveguide Crossing" sch_x=54 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C553 N$2064 N$2066 N$2017 N$2019 "Waveguide Crossing" sch_x=54 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C554 N$2068 N$2070 N$2021 N$2023 "Waveguide Crossing" sch_x=54 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C555 N$2072 N$2074 N$2025 N$2027 "Waveguide Crossing" sch_x=54 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C556 N$2076 N$2078 N$2029 N$2031 "Waveguide Crossing" sch_x=54 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C557 N$2080 N$2082 N$2033 N$2035 "Waveguide Crossing" sch_x=54 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C558 N$2084 N$2357 N$2037 N$2039 "Waveguide Crossing" sch_x=54 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C559 N$2313 N$2086 N$2041 N$2043 "Waveguide Crossing" sch_x=52 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C560 N$2088 N$2090 N$2045 N$2047 "Waveguide Crossing" sch_x=52 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C561 N$2092 N$2094 N$2049 N$2051 "Waveguide Crossing" sch_x=52 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C562 N$2096 N$2098 N$2053 N$2055 "Waveguide Crossing" sch_x=52 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C563 N$2100 N$2102 N$2057 N$2059 "Waveguide Crossing" sch_x=52 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C564 N$2104 N$2106 N$2061 N$2063 "Waveguide Crossing" sch_x=52 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C565 N$2108 N$2110 N$2065 N$2067 "Waveguide Crossing" sch_x=52 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C566 N$2112 N$2114 N$2069 N$2071 "Waveguide Crossing" sch_x=52 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C567 N$2116 N$2118 N$2073 N$2075 "Waveguide Crossing" sch_x=52 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C568 N$2120 N$2122 N$2077 N$2079 "Waveguide Crossing" sch_x=52 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C569 N$2124 N$2355 N$2081 N$2083 "Waveguide Crossing" sch_x=52 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C570 N$2315 N$2126 N$2085 N$2087 "Waveguide Crossing" sch_x=50 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C571 N$2128 N$2130 N$2089 N$2091 "Waveguide Crossing" sch_x=50 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C572 N$2132 N$2134 N$2093 N$2095 "Waveguide Crossing" sch_x=50 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C573 N$2136 N$2138 N$2097 N$2099 "Waveguide Crossing" sch_x=50 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C574 N$2140 N$2142 N$2101 N$2103 "Waveguide Crossing" sch_x=50 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C575 N$2144 N$2146 N$2105 N$2107 "Waveguide Crossing" sch_x=50 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C576 N$2148 N$2150 N$2109 N$2111 "Waveguide Crossing" sch_x=50 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C577 N$2152 N$2154 N$2113 N$2115 "Waveguide Crossing" sch_x=50 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C578 N$2156 N$2158 N$2117 N$2119 "Waveguide Crossing" sch_x=50 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C579 N$2160 N$2353 N$2121 N$2123 "Waveguide Crossing" sch_x=50 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C580 N$2317 N$2162 N$2125 N$2127 "Waveguide Crossing" sch_x=48 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C581 N$2164 N$2166 N$2129 N$2131 "Waveguide Crossing" sch_x=48 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C582 N$2168 N$2170 N$2133 N$2135 "Waveguide Crossing" sch_x=48 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C583 N$2172 N$2174 N$2137 N$2139 "Waveguide Crossing" sch_x=48 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C584 N$2176 N$2178 N$2141 N$2143 "Waveguide Crossing" sch_x=48 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C585 N$2180 N$2182 N$2145 N$2147 "Waveguide Crossing" sch_x=48 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C586 N$2184 N$2186 N$2149 N$2151 "Waveguide Crossing" sch_x=48 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C587 N$2188 N$2190 N$2153 N$2155 "Waveguide Crossing" sch_x=48 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C588 N$2192 N$2351 N$2157 N$2159 "Waveguide Crossing" sch_x=48 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C589 N$2319 N$2194 N$2161 N$2163 "Waveguide Crossing" sch_x=46 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C590 N$2196 N$2198 N$2165 N$2167 "Waveguide Crossing" sch_x=46 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C591 N$2200 N$2202 N$2169 N$2171 "Waveguide Crossing" sch_x=46 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C592 N$2204 N$2206 N$2173 N$2175 "Waveguide Crossing" sch_x=46 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C593 N$2208 N$2210 N$2177 N$2179 "Waveguide Crossing" sch_x=46 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C594 N$2212 N$2214 N$2181 N$2183 "Waveguide Crossing" sch_x=46 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C595 N$2216 N$2218 N$2185 N$2187 "Waveguide Crossing" sch_x=46 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C596 N$2220 N$2349 N$2189 N$2191 "Waveguide Crossing" sch_x=46 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C597 N$2321 N$2222 N$2193 N$2195 "Waveguide Crossing" sch_x=44 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C598 N$2224 N$2226 N$2197 N$2199 "Waveguide Crossing" sch_x=44 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C599 N$2228 N$2230 N$2201 N$2203 "Waveguide Crossing" sch_x=44 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C600 N$2232 N$2234 N$2205 N$2207 "Waveguide Crossing" sch_x=44 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C601 N$2236 N$2238 N$2209 N$2211 "Waveguide Crossing" sch_x=44 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C602 N$2240 N$2242 N$2213 N$2215 "Waveguide Crossing" sch_x=44 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C603 N$2244 N$2347 N$2217 N$2219 "Waveguide Crossing" sch_x=44 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C604 N$2323 N$2246 N$2221 N$2223 "Waveguide Crossing" sch_x=42 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C605 N$2248 N$2250 N$2225 N$2227 "Waveguide Crossing" sch_x=42 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C606 N$2252 N$2254 N$2229 N$2231 "Waveguide Crossing" sch_x=42 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C607 N$2256 N$2258 N$2233 N$2235 "Waveguide Crossing" sch_x=42 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C608 N$2260 N$2262 N$2237 N$2239 "Waveguide Crossing" sch_x=42 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C609 N$2264 N$2345 N$2241 N$2243 "Waveguide Crossing" sch_x=42 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C610 N$2325 N$2266 N$2245 N$2247 "Waveguide Crossing" sch_x=40 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C611 N$2268 N$2270 N$2249 N$2251 "Waveguide Crossing" sch_x=40 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C612 N$2272 N$2274 N$2253 N$2255 "Waveguide Crossing" sch_x=40 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C613 N$2276 N$2278 N$2257 N$2259 "Waveguide Crossing" sch_x=40 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C614 N$2280 N$2343 N$2261 N$2263 "Waveguide Crossing" sch_x=40 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C615 N$2327 N$2282 N$2265 N$2267 "Waveguide Crossing" sch_x=38 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C616 N$2284 N$2286 N$2269 N$2271 "Waveguide Crossing" sch_x=38 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C617 N$2288 N$2290 N$2273 N$2275 "Waveguide Crossing" sch_x=38 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C618 N$2292 N$2341 N$2277 N$2279 "Waveguide Crossing" sch_x=38 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C619 N$2329 N$2294 N$2281 N$2283 "Waveguide Crossing" sch_x=36 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C620 N$2296 N$2298 N$2285 N$2287 "Waveguide Crossing" sch_x=36 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C621 N$2300 N$2339 N$2289 N$2291 "Waveguide Crossing" sch_x=36 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C622 N$2331 N$2302 N$2293 N$2295 "Waveguide Crossing" sch_x=34 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C623 N$2304 N$2337 N$2297 N$2299 "Waveguide Crossing" sch_x=34 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C624 N$2333 N$2335 N$2301 N$2303 "Waveguide Crossing" sch_x=32 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S489 N$2365 N$1826 N$8958 N$8834 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S490 N$1828 N$1830 N$8836 N$8838 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S491 N$1832 N$1834 N$8840 N$8842 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S492 N$1836 N$1838 N$8844 N$8846 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S493 N$1840 N$1842 N$8848 N$8850 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S494 N$1844 N$1846 N$8852 N$8854 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S495 N$1848 N$1850 N$8856 N$8858 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S496 N$1852 N$1854 N$8860 N$8862 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S497 N$1856 N$1858 N$8864 N$8866 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S498 N$1860 N$1862 N$8868 N$8870 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S499 N$1864 N$1866 N$8872 N$8874 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S500 N$1868 N$1870 N$8876 N$8878 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S501 N$1872 N$1874 N$8880 N$8882 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S502 N$1876 N$1878 N$8884 N$8886 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S503 N$1880 N$1882 N$8888 N$8890 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S504 N$1884 N$2367 N$8892 N$8894 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S625 N$2502 N$2490 N$2369 N$2371 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S626 N$2492 N$2494 N$2373 N$2379 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S627 N$34753 N$2370 N$2381 N$2383 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S628 N$2376 N$34754 N$2385 N$2391 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S629 N$34755 N$2378 N$2393 N$2395 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S630 N$2380 N$34756 N$2397 N$2403 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S631 N$2382 N$2390 N$2405 N$34757 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S632 N$2388 N$2392 N$34758 N$2407 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S633 N$2394 N$2402 N$2409 N$34759 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S634 N$2400 N$2404 N$34760 N$2415 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S635 N$2406 N$2414 N$2542 N$2530 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S636 N$2412 N$2416 N$2532 N$2534 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C637 N$2372 N$2374 N$2375 N$2377 "Waveguide Crossing" sch_x=-4 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C638 N$2384 N$2386 N$2389 N$2387 "Waveguide Crossing" sch_x=0 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C639 N$2396 N$2398 N$2401 N$2399 "Waveguide Crossing" sch_x=0 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C640 N$2408 N$2410 N$2413 N$2411 "Waveguide Crossing" sch_x=4 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S641 N$2496 N$2498 N$2417 N$2419 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S642 N$2500 N$2504 N$2421 N$2427 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S643 N$34761 N$2418 N$2429 N$2431 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S644 N$2424 N$34762 N$2433 N$2439 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S645 N$34763 N$2426 N$2441 N$2443 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S646 N$2428 N$34764 N$2445 N$2451 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S647 N$2430 N$2438 N$2453 N$34765 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S648 N$2436 N$2440 N$34766 N$2455 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S649 N$2442 N$2450 N$2457 N$34767 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S650 N$2448 N$2452 N$34768 N$2463 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S651 N$2454 N$2462 N$2536 N$2538 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S652 N$2460 N$2464 N$2540 N$2544 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C653 N$2420 N$2422 N$2423 N$2425 "Waveguide Crossing" sch_x=-4 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C654 N$2432 N$2434 N$2437 N$2435 "Waveguide Crossing" sch_x=0 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C655 N$2444 N$2446 N$2449 N$2447 "Waveguide Crossing" sch_x=0 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C656 N$2456 N$2458 N$2461 N$2459 "Waveguide Crossing" sch_x=4 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C671 N$2529 N$2518 N$2505 N$2507 "Waveguide Crossing" sch_x=12 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C672 N$2520 N$2522 N$2509 N$2511 "Waveguide Crossing" sch_x=12 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C673 N$2524 N$2539 N$2513 N$2515 "Waveguide Crossing" sch_x=12 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C674 N$2531 N$2526 N$2517 N$2519 "Waveguide Crossing" sch_x=10 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C675 N$2528 N$2537 N$2521 N$2523 "Waveguide Crossing" sch_x=10 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C676 N$2533 N$2535 N$2525 N$2527 "Waveguide Crossing" sch_x=8 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S667 N$2541 N$2506 N$3006 N$2978 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S668 N$2508 N$2510 N$2980 N$2982 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S669 N$2512 N$2514 N$2984 N$2986 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S670 N$2516 N$2543 N$2988 N$2990 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S677 N$2678 N$2666 N$2545 N$2547 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S678 N$2668 N$2670 N$2549 N$2555 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S679 N$34769 N$2546 N$2557 N$2559 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S680 N$2552 N$34770 N$2561 N$2567 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S681 N$34771 N$2554 N$2569 N$2571 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S682 N$2556 N$34772 N$2573 N$2579 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S683 N$2558 N$2566 N$2581 N$34773 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S684 N$2564 N$2568 N$34774 N$2583 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S685 N$2570 N$2578 N$2585 N$34775 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S686 N$2576 N$2580 N$34776 N$2591 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S687 N$2582 N$2590 N$2718 N$2706 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S688 N$2588 N$2592 N$2708 N$2710 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C689 N$2548 N$2550 N$2551 N$2553 "Waveguide Crossing" sch_x=-4 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C690 N$2560 N$2562 N$2565 N$2563 "Waveguide Crossing" sch_x=0 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C691 N$2572 N$2574 N$2577 N$2575 "Waveguide Crossing" sch_x=0 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C692 N$2584 N$2586 N$2589 N$2587 "Waveguide Crossing" sch_x=4 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S693 N$2672 N$2674 N$2593 N$2595 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S694 N$2676 N$2680 N$2597 N$2603 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S695 N$34777 N$2594 N$2605 N$2607 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S696 N$2600 N$34778 N$2609 N$2615 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S697 N$34779 N$2602 N$2617 N$2619 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S698 N$2604 N$34780 N$2621 N$2627 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S699 N$2606 N$2614 N$2629 N$34781 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S700 N$2612 N$2616 N$34782 N$2631 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S701 N$2618 N$2626 N$2633 N$34783 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S702 N$2624 N$2628 N$34784 N$2639 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S703 N$2630 N$2638 N$2712 N$2714 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S704 N$2636 N$2640 N$2716 N$2720 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C705 N$2596 N$2598 N$2599 N$2601 "Waveguide Crossing" sch_x=-4 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C706 N$2608 N$2610 N$2613 N$2611 "Waveguide Crossing" sch_x=0 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C707 N$2620 N$2622 N$2625 N$2623 "Waveguide Crossing" sch_x=0 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C708 N$2632 N$2634 N$2637 N$2635 "Waveguide Crossing" sch_x=4 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C723 N$2705 N$2694 N$2681 N$2683 "Waveguide Crossing" sch_x=12 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C724 N$2696 N$2698 N$2685 N$2687 "Waveguide Crossing" sch_x=12 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C725 N$2700 N$2715 N$2689 N$2691 "Waveguide Crossing" sch_x=12 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C726 N$2707 N$2702 N$2693 N$2695 "Waveguide Crossing" sch_x=10 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C727 N$2704 N$2713 N$2697 N$2699 "Waveguide Crossing" sch_x=10 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C728 N$2709 N$2711 N$2701 N$2703 "Waveguide Crossing" sch_x=8 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S719 N$2717 N$2682 N$2992 N$2994 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S720 N$2684 N$2686 N$2996 N$2998 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S721 N$2688 N$2690 N$3000 N$3002 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S722 N$2692 N$2719 N$3004 N$3008 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C773 N$2977 N$2894 N$2865 N$2867 "Waveguide Crossing" sch_x=28 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C774 N$2896 N$2898 N$2869 N$2871 "Waveguide Crossing" sch_x=28 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C775 N$2900 N$2902 N$2873 N$2875 "Waveguide Crossing" sch_x=28 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C776 N$2904 N$2906 N$2877 N$2879 "Waveguide Crossing" sch_x=28 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C777 N$2908 N$2910 N$2881 N$2883 "Waveguide Crossing" sch_x=28 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C778 N$2912 N$2914 N$2885 N$2887 "Waveguide Crossing" sch_x=28 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C779 N$2916 N$3003 N$2889 N$2891 "Waveguide Crossing" sch_x=28 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C780 N$2979 N$2918 N$2893 N$2895 "Waveguide Crossing" sch_x=26 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C781 N$2920 N$2922 N$2897 N$2899 "Waveguide Crossing" sch_x=26 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C782 N$2924 N$2926 N$2901 N$2903 "Waveguide Crossing" sch_x=26 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C783 N$2928 N$2930 N$2905 N$2907 "Waveguide Crossing" sch_x=26 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C784 N$2932 N$2934 N$2909 N$2911 "Waveguide Crossing" sch_x=26 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C785 N$2936 N$3001 N$2913 N$2915 "Waveguide Crossing" sch_x=26 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C786 N$2981 N$2938 N$2917 N$2919 "Waveguide Crossing" sch_x=24 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C787 N$2940 N$2942 N$2921 N$2923 "Waveguide Crossing" sch_x=24 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C788 N$2944 N$2946 N$2925 N$2927 "Waveguide Crossing" sch_x=24 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C789 N$2948 N$2950 N$2929 N$2931 "Waveguide Crossing" sch_x=24 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C790 N$2952 N$2999 N$2933 N$2935 "Waveguide Crossing" sch_x=24 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C791 N$2983 N$2954 N$2937 N$2939 "Waveguide Crossing" sch_x=22 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C792 N$2956 N$2958 N$2941 N$2943 "Waveguide Crossing" sch_x=22 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C793 N$2960 N$2962 N$2945 N$2947 "Waveguide Crossing" sch_x=22 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C794 N$2964 N$2997 N$2949 N$2951 "Waveguide Crossing" sch_x=22 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C795 N$2985 N$2966 N$2953 N$2955 "Waveguide Crossing" sch_x=20 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C796 N$2968 N$2970 N$2957 N$2959 "Waveguide Crossing" sch_x=20 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C797 N$2972 N$2995 N$2961 N$2963 "Waveguide Crossing" sch_x=20 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C798 N$2987 N$2974 N$2965 N$2967 "Waveguide Crossing" sch_x=18 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C799 N$2976 N$2993 N$2969 N$2971 "Waveguide Crossing" sch_x=18 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C800 N$2989 N$2991 N$2973 N$2975 "Waveguide Crossing" sch_x=16 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S765 N$3005 N$2866 N$4734 N$4674 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S766 N$2868 N$2870 N$4676 N$4678 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S767 N$2872 N$2874 N$4680 N$4682 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S768 N$2876 N$2878 N$4684 N$4686 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S769 N$2880 N$2882 N$4688 N$4690 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S770 N$2884 N$2886 N$4692 N$4694 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S771 N$2888 N$2890 N$4696 N$4698 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S772 N$2892 N$3007 N$4700 N$4702 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S801 N$3142 N$3130 N$3009 N$3011 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S802 N$3132 N$3134 N$3013 N$3019 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S803 N$34785 N$3010 N$3021 N$3023 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S804 N$3016 N$34786 N$3025 N$3031 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S805 N$34787 N$3018 N$3033 N$3035 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S806 N$3020 N$34788 N$3037 N$3043 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S807 N$3022 N$3030 N$3045 N$34789 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S808 N$3028 N$3032 N$34790 N$3047 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S809 N$3034 N$3042 N$3049 N$34791 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S810 N$3040 N$3044 N$34792 N$3055 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S811 N$3046 N$3054 N$3182 N$3170 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S812 N$3052 N$3056 N$3172 N$3174 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C813 N$3012 N$3014 N$3015 N$3017 "Waveguide Crossing" sch_x=-4 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C814 N$3024 N$3026 N$3029 N$3027 "Waveguide Crossing" sch_x=0 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C815 N$3036 N$3038 N$3041 N$3039 "Waveguide Crossing" sch_x=0 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C816 N$3048 N$3050 N$3053 N$3051 "Waveguide Crossing" sch_x=4 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S817 N$3136 N$3138 N$3057 N$3059 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S818 N$3140 N$3144 N$3061 N$3067 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S819 N$34793 N$3058 N$3069 N$3071 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S820 N$3064 N$34794 N$3073 N$3079 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S821 N$34795 N$3066 N$3081 N$3083 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S822 N$3068 N$34796 N$3085 N$3091 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S823 N$3070 N$3078 N$3093 N$34797 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S824 N$3076 N$3080 N$34798 N$3095 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S825 N$3082 N$3090 N$3097 N$34799 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S826 N$3088 N$3092 N$34800 N$3103 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S827 N$3094 N$3102 N$3176 N$3178 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S828 N$3100 N$3104 N$3180 N$3184 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C829 N$3060 N$3062 N$3063 N$3065 "Waveguide Crossing" sch_x=-4 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C830 N$3072 N$3074 N$3077 N$3075 "Waveguide Crossing" sch_x=0 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C831 N$3084 N$3086 N$3089 N$3087 "Waveguide Crossing" sch_x=0 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C832 N$3096 N$3098 N$3101 N$3099 "Waveguide Crossing" sch_x=4 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C847 N$3169 N$3158 N$3145 N$3147 "Waveguide Crossing" sch_x=12 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C848 N$3160 N$3162 N$3149 N$3151 "Waveguide Crossing" sch_x=12 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C849 N$3164 N$3179 N$3153 N$3155 "Waveguide Crossing" sch_x=12 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C850 N$3171 N$3166 N$3157 N$3159 "Waveguide Crossing" sch_x=10 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C851 N$3168 N$3177 N$3161 N$3163 "Waveguide Crossing" sch_x=10 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C852 N$3173 N$3175 N$3165 N$3167 "Waveguide Crossing" sch_x=8 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S843 N$3181 N$3146 N$3646 N$3618 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S844 N$3148 N$3150 N$3620 N$3622 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S845 N$3152 N$3154 N$3624 N$3626 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S846 N$3156 N$3183 N$3628 N$3630 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S853 N$3318 N$3306 N$3185 N$3187 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S854 N$3308 N$3310 N$3189 N$3195 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S855 N$34801 N$3186 N$3197 N$3199 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S856 N$3192 N$34802 N$3201 N$3207 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S857 N$34803 N$3194 N$3209 N$3211 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S858 N$3196 N$34804 N$3213 N$3219 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S859 N$3198 N$3206 N$3221 N$34805 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S860 N$3204 N$3208 N$34806 N$3223 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S861 N$3210 N$3218 N$3225 N$34807 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S862 N$3216 N$3220 N$34808 N$3231 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S863 N$3222 N$3230 N$3358 N$3346 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S864 N$3228 N$3232 N$3348 N$3350 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C865 N$3188 N$3190 N$3191 N$3193 "Waveguide Crossing" sch_x=-4 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C866 N$3200 N$3202 N$3205 N$3203 "Waveguide Crossing" sch_x=0 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C867 N$3212 N$3214 N$3217 N$3215 "Waveguide Crossing" sch_x=0 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C868 N$3224 N$3226 N$3229 N$3227 "Waveguide Crossing" sch_x=4 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S869 N$3312 N$3314 N$3233 N$3235 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S870 N$3316 N$3320 N$3237 N$3243 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S871 N$34809 N$3234 N$3245 N$3247 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S872 N$3240 N$34810 N$3249 N$3255 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S873 N$34811 N$3242 N$3257 N$3259 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S874 N$3244 N$34812 N$3261 N$3267 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S875 N$3246 N$3254 N$3269 N$34813 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S876 N$3252 N$3256 N$34814 N$3271 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S877 N$3258 N$3266 N$3273 N$34815 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S878 N$3264 N$3268 N$34816 N$3279 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S879 N$3270 N$3278 N$3352 N$3354 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S880 N$3276 N$3280 N$3356 N$3360 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C881 N$3236 N$3238 N$3239 N$3241 "Waveguide Crossing" sch_x=-4 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C882 N$3248 N$3250 N$3253 N$3251 "Waveguide Crossing" sch_x=0 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C883 N$3260 N$3262 N$3265 N$3263 "Waveguide Crossing" sch_x=0 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C884 N$3272 N$3274 N$3277 N$3275 "Waveguide Crossing" sch_x=4 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C899 N$3345 N$3334 N$3321 N$3323 "Waveguide Crossing" sch_x=12 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C900 N$3336 N$3338 N$3325 N$3327 "Waveguide Crossing" sch_x=12 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C901 N$3340 N$3355 N$3329 N$3331 "Waveguide Crossing" sch_x=12 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C902 N$3347 N$3342 N$3333 N$3335 "Waveguide Crossing" sch_x=10 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C903 N$3344 N$3353 N$3337 N$3339 "Waveguide Crossing" sch_x=10 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C904 N$3349 N$3351 N$3341 N$3343 "Waveguide Crossing" sch_x=8 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S895 N$3357 N$3322 N$3632 N$3634 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S896 N$3324 N$3326 N$3636 N$3638 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S897 N$3328 N$3330 N$3640 N$3642 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S898 N$3332 N$3359 N$3644 N$3648 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C949 N$3617 N$3534 N$3505 N$3507 "Waveguide Crossing" sch_x=28 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C950 N$3536 N$3538 N$3509 N$3511 "Waveguide Crossing" sch_x=28 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C951 N$3540 N$3542 N$3513 N$3515 "Waveguide Crossing" sch_x=28 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C952 N$3544 N$3546 N$3517 N$3519 "Waveguide Crossing" sch_x=28 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C953 N$3548 N$3550 N$3521 N$3523 "Waveguide Crossing" sch_x=28 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C954 N$3552 N$3554 N$3525 N$3527 "Waveguide Crossing" sch_x=28 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C955 N$3556 N$3643 N$3529 N$3531 "Waveguide Crossing" sch_x=28 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C956 N$3619 N$3558 N$3533 N$3535 "Waveguide Crossing" sch_x=26 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C957 N$3560 N$3562 N$3537 N$3539 "Waveguide Crossing" sch_x=26 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C958 N$3564 N$3566 N$3541 N$3543 "Waveguide Crossing" sch_x=26 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C959 N$3568 N$3570 N$3545 N$3547 "Waveguide Crossing" sch_x=26 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C960 N$3572 N$3574 N$3549 N$3551 "Waveguide Crossing" sch_x=26 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C961 N$3576 N$3641 N$3553 N$3555 "Waveguide Crossing" sch_x=26 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C962 N$3621 N$3578 N$3557 N$3559 "Waveguide Crossing" sch_x=24 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C963 N$3580 N$3582 N$3561 N$3563 "Waveguide Crossing" sch_x=24 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C964 N$3584 N$3586 N$3565 N$3567 "Waveguide Crossing" sch_x=24 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C965 N$3588 N$3590 N$3569 N$3571 "Waveguide Crossing" sch_x=24 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C966 N$3592 N$3639 N$3573 N$3575 "Waveguide Crossing" sch_x=24 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C967 N$3623 N$3594 N$3577 N$3579 "Waveguide Crossing" sch_x=22 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C968 N$3596 N$3598 N$3581 N$3583 "Waveguide Crossing" sch_x=22 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C969 N$3600 N$3602 N$3585 N$3587 "Waveguide Crossing" sch_x=22 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C970 N$3604 N$3637 N$3589 N$3591 "Waveguide Crossing" sch_x=22 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C971 N$3625 N$3606 N$3593 N$3595 "Waveguide Crossing" sch_x=20 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C972 N$3608 N$3610 N$3597 N$3599 "Waveguide Crossing" sch_x=20 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C973 N$3612 N$3635 N$3601 N$3603 "Waveguide Crossing" sch_x=20 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C974 N$3627 N$3614 N$3605 N$3607 "Waveguide Crossing" sch_x=18 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C975 N$3616 N$3633 N$3609 N$3611 "Waveguide Crossing" sch_x=18 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C976 N$3629 N$3631 N$3613 N$3615 "Waveguide Crossing" sch_x=16 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S941 N$3645 N$3506 N$4704 N$4706 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S942 N$3508 N$3510 N$4708 N$4710 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S943 N$3512 N$3514 N$4712 N$4714 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S944 N$3516 N$3518 N$4716 N$4718 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S945 N$3520 N$3522 N$4720 N$4722 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S946 N$3524 N$3526 N$4724 N$4726 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S947 N$3528 N$3530 N$4728 N$4730 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S948 N$3532 N$3647 N$4732 N$4736 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1129 N$4673 N$4254 N$4193 N$4195 "Waveguide Crossing" sch_x=60 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1130 N$4256 N$4258 N$4197 N$4199 "Waveguide Crossing" sch_x=60 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1131 N$4260 N$4262 N$4201 N$4203 "Waveguide Crossing" sch_x=60 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1132 N$4264 N$4266 N$4205 N$4207 "Waveguide Crossing" sch_x=60 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1133 N$4268 N$4270 N$4209 N$4211 "Waveguide Crossing" sch_x=60 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1134 N$4272 N$4274 N$4213 N$4215 "Waveguide Crossing" sch_x=60 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1135 N$4276 N$4278 N$4217 N$4219 "Waveguide Crossing" sch_x=60 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1136 N$4280 N$4282 N$4221 N$4223 "Waveguide Crossing" sch_x=60 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1137 N$4284 N$4286 N$4225 N$4227 "Waveguide Crossing" sch_x=60 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1138 N$4288 N$4290 N$4229 N$4231 "Waveguide Crossing" sch_x=60 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1139 N$4292 N$4294 N$4233 N$4235 "Waveguide Crossing" sch_x=60 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1140 N$4296 N$4298 N$4237 N$4239 "Waveguide Crossing" sch_x=60 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1141 N$4300 N$4302 N$4241 N$4243 "Waveguide Crossing" sch_x=60 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1142 N$4304 N$4306 N$4245 N$4247 "Waveguide Crossing" sch_x=60 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1143 N$4308 N$4731 N$4249 N$4251 "Waveguide Crossing" sch_x=60 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1144 N$4675 N$4310 N$4253 N$4255 "Waveguide Crossing" sch_x=58 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1145 N$4312 N$4314 N$4257 N$4259 "Waveguide Crossing" sch_x=58 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1146 N$4316 N$4318 N$4261 N$4263 "Waveguide Crossing" sch_x=58 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1147 N$4320 N$4322 N$4265 N$4267 "Waveguide Crossing" sch_x=58 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1148 N$4324 N$4326 N$4269 N$4271 "Waveguide Crossing" sch_x=58 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1149 N$4328 N$4330 N$4273 N$4275 "Waveguide Crossing" sch_x=58 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1150 N$4332 N$4334 N$4277 N$4279 "Waveguide Crossing" sch_x=58 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1151 N$4336 N$4338 N$4281 N$4283 "Waveguide Crossing" sch_x=58 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1152 N$4340 N$4342 N$4285 N$4287 "Waveguide Crossing" sch_x=58 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1153 N$4344 N$4346 N$4289 N$4291 "Waveguide Crossing" sch_x=58 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1154 N$4348 N$4350 N$4293 N$4295 "Waveguide Crossing" sch_x=58 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1155 N$4352 N$4354 N$4297 N$4299 "Waveguide Crossing" sch_x=58 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1156 N$4356 N$4358 N$4301 N$4303 "Waveguide Crossing" sch_x=58 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1157 N$4360 N$4729 N$4305 N$4307 "Waveguide Crossing" sch_x=58 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1158 N$4677 N$4362 N$4309 N$4311 "Waveguide Crossing" sch_x=56 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1159 N$4364 N$4366 N$4313 N$4315 "Waveguide Crossing" sch_x=56 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1160 N$4368 N$4370 N$4317 N$4319 "Waveguide Crossing" sch_x=56 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1161 N$4372 N$4374 N$4321 N$4323 "Waveguide Crossing" sch_x=56 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1162 N$4376 N$4378 N$4325 N$4327 "Waveguide Crossing" sch_x=56 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1163 N$4380 N$4382 N$4329 N$4331 "Waveguide Crossing" sch_x=56 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1164 N$4384 N$4386 N$4333 N$4335 "Waveguide Crossing" sch_x=56 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1165 N$4388 N$4390 N$4337 N$4339 "Waveguide Crossing" sch_x=56 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1166 N$4392 N$4394 N$4341 N$4343 "Waveguide Crossing" sch_x=56 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1167 N$4396 N$4398 N$4345 N$4347 "Waveguide Crossing" sch_x=56 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1168 N$4400 N$4402 N$4349 N$4351 "Waveguide Crossing" sch_x=56 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1169 N$4404 N$4406 N$4353 N$4355 "Waveguide Crossing" sch_x=56 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1170 N$4408 N$4727 N$4357 N$4359 "Waveguide Crossing" sch_x=56 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1171 N$4679 N$4410 N$4361 N$4363 "Waveguide Crossing" sch_x=54 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1172 N$4412 N$4414 N$4365 N$4367 "Waveguide Crossing" sch_x=54 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1173 N$4416 N$4418 N$4369 N$4371 "Waveguide Crossing" sch_x=54 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1174 N$4420 N$4422 N$4373 N$4375 "Waveguide Crossing" sch_x=54 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1175 N$4424 N$4426 N$4377 N$4379 "Waveguide Crossing" sch_x=54 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1176 N$4428 N$4430 N$4381 N$4383 "Waveguide Crossing" sch_x=54 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1177 N$4432 N$4434 N$4385 N$4387 "Waveguide Crossing" sch_x=54 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1178 N$4436 N$4438 N$4389 N$4391 "Waveguide Crossing" sch_x=54 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1179 N$4440 N$4442 N$4393 N$4395 "Waveguide Crossing" sch_x=54 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1180 N$4444 N$4446 N$4397 N$4399 "Waveguide Crossing" sch_x=54 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1181 N$4448 N$4450 N$4401 N$4403 "Waveguide Crossing" sch_x=54 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1182 N$4452 N$4725 N$4405 N$4407 "Waveguide Crossing" sch_x=54 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1183 N$4681 N$4454 N$4409 N$4411 "Waveguide Crossing" sch_x=52 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1184 N$4456 N$4458 N$4413 N$4415 "Waveguide Crossing" sch_x=52 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1185 N$4460 N$4462 N$4417 N$4419 "Waveguide Crossing" sch_x=52 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1186 N$4464 N$4466 N$4421 N$4423 "Waveguide Crossing" sch_x=52 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1187 N$4468 N$4470 N$4425 N$4427 "Waveguide Crossing" sch_x=52 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1188 N$4472 N$4474 N$4429 N$4431 "Waveguide Crossing" sch_x=52 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1189 N$4476 N$4478 N$4433 N$4435 "Waveguide Crossing" sch_x=52 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1190 N$4480 N$4482 N$4437 N$4439 "Waveguide Crossing" sch_x=52 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1191 N$4484 N$4486 N$4441 N$4443 "Waveguide Crossing" sch_x=52 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1192 N$4488 N$4490 N$4445 N$4447 "Waveguide Crossing" sch_x=52 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1193 N$4492 N$4723 N$4449 N$4451 "Waveguide Crossing" sch_x=52 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1194 N$4683 N$4494 N$4453 N$4455 "Waveguide Crossing" sch_x=50 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1195 N$4496 N$4498 N$4457 N$4459 "Waveguide Crossing" sch_x=50 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1196 N$4500 N$4502 N$4461 N$4463 "Waveguide Crossing" sch_x=50 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1197 N$4504 N$4506 N$4465 N$4467 "Waveguide Crossing" sch_x=50 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1198 N$4508 N$4510 N$4469 N$4471 "Waveguide Crossing" sch_x=50 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1199 N$4512 N$4514 N$4473 N$4475 "Waveguide Crossing" sch_x=50 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1200 N$4516 N$4518 N$4477 N$4479 "Waveguide Crossing" sch_x=50 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1201 N$4520 N$4522 N$4481 N$4483 "Waveguide Crossing" sch_x=50 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1202 N$4524 N$4526 N$4485 N$4487 "Waveguide Crossing" sch_x=50 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1203 N$4528 N$4721 N$4489 N$4491 "Waveguide Crossing" sch_x=50 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1204 N$4685 N$4530 N$4493 N$4495 "Waveguide Crossing" sch_x=48 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1205 N$4532 N$4534 N$4497 N$4499 "Waveguide Crossing" sch_x=48 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1206 N$4536 N$4538 N$4501 N$4503 "Waveguide Crossing" sch_x=48 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1207 N$4540 N$4542 N$4505 N$4507 "Waveguide Crossing" sch_x=48 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1208 N$4544 N$4546 N$4509 N$4511 "Waveguide Crossing" sch_x=48 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1209 N$4548 N$4550 N$4513 N$4515 "Waveguide Crossing" sch_x=48 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1210 N$4552 N$4554 N$4517 N$4519 "Waveguide Crossing" sch_x=48 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1211 N$4556 N$4558 N$4521 N$4523 "Waveguide Crossing" sch_x=48 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1212 N$4560 N$4719 N$4525 N$4527 "Waveguide Crossing" sch_x=48 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1213 N$4687 N$4562 N$4529 N$4531 "Waveguide Crossing" sch_x=46 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1214 N$4564 N$4566 N$4533 N$4535 "Waveguide Crossing" sch_x=46 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1215 N$4568 N$4570 N$4537 N$4539 "Waveguide Crossing" sch_x=46 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1216 N$4572 N$4574 N$4541 N$4543 "Waveguide Crossing" sch_x=46 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1217 N$4576 N$4578 N$4545 N$4547 "Waveguide Crossing" sch_x=46 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1218 N$4580 N$4582 N$4549 N$4551 "Waveguide Crossing" sch_x=46 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1219 N$4584 N$4586 N$4553 N$4555 "Waveguide Crossing" sch_x=46 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1220 N$4588 N$4717 N$4557 N$4559 "Waveguide Crossing" sch_x=46 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1221 N$4689 N$4590 N$4561 N$4563 "Waveguide Crossing" sch_x=44 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1222 N$4592 N$4594 N$4565 N$4567 "Waveguide Crossing" sch_x=44 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1223 N$4596 N$4598 N$4569 N$4571 "Waveguide Crossing" sch_x=44 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1224 N$4600 N$4602 N$4573 N$4575 "Waveguide Crossing" sch_x=44 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1225 N$4604 N$4606 N$4577 N$4579 "Waveguide Crossing" sch_x=44 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1226 N$4608 N$4610 N$4581 N$4583 "Waveguide Crossing" sch_x=44 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1227 N$4612 N$4715 N$4585 N$4587 "Waveguide Crossing" sch_x=44 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1228 N$4691 N$4614 N$4589 N$4591 "Waveguide Crossing" sch_x=42 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1229 N$4616 N$4618 N$4593 N$4595 "Waveguide Crossing" sch_x=42 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1230 N$4620 N$4622 N$4597 N$4599 "Waveguide Crossing" sch_x=42 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1231 N$4624 N$4626 N$4601 N$4603 "Waveguide Crossing" sch_x=42 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1232 N$4628 N$4630 N$4605 N$4607 "Waveguide Crossing" sch_x=42 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1233 N$4632 N$4713 N$4609 N$4611 "Waveguide Crossing" sch_x=42 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1234 N$4693 N$4634 N$4613 N$4615 "Waveguide Crossing" sch_x=40 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1235 N$4636 N$4638 N$4617 N$4619 "Waveguide Crossing" sch_x=40 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1236 N$4640 N$4642 N$4621 N$4623 "Waveguide Crossing" sch_x=40 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1237 N$4644 N$4646 N$4625 N$4627 "Waveguide Crossing" sch_x=40 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1238 N$4648 N$4711 N$4629 N$4631 "Waveguide Crossing" sch_x=40 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1239 N$4695 N$4650 N$4633 N$4635 "Waveguide Crossing" sch_x=38 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1240 N$4652 N$4654 N$4637 N$4639 "Waveguide Crossing" sch_x=38 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1241 N$4656 N$4658 N$4641 N$4643 "Waveguide Crossing" sch_x=38 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1242 N$4660 N$4709 N$4645 N$4647 "Waveguide Crossing" sch_x=38 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1243 N$4697 N$4662 N$4649 N$4651 "Waveguide Crossing" sch_x=36 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1244 N$4664 N$4666 N$4653 N$4655 "Waveguide Crossing" sch_x=36 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1245 N$4668 N$4707 N$4657 N$4659 "Waveguide Crossing" sch_x=36 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1246 N$4699 N$4670 N$4661 N$4663 "Waveguide Crossing" sch_x=34 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1247 N$4672 N$4705 N$4665 N$4667 "Waveguide Crossing" sch_x=34 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1248 N$4701 N$4703 N$4669 N$4671 "Waveguide Crossing" sch_x=32 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1113 N$4733 N$4194 N$8896 N$8898 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1114 N$4196 N$4198 N$8900 N$8902 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1115 N$4200 N$4202 N$8904 N$8906 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1116 N$4204 N$4206 N$8908 N$8910 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1117 N$4208 N$4210 N$8912 N$8914 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1118 N$4212 N$4214 N$8916 N$8918 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1119 N$4216 N$4218 N$8920 N$8922 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1120 N$4220 N$4222 N$8924 N$8926 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1121 N$4224 N$4226 N$8928 N$8930 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1122 N$4228 N$4230 N$8932 N$8934 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1123 N$4232 N$4234 N$8936 N$8938 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1124 N$4236 N$4238 N$8940 N$8942 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1125 N$4240 N$4242 N$8944 N$8946 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1126 N$4244 N$4246 N$8948 N$8950 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1127 N$4248 N$4250 N$8952 N$8954 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1128 N$4252 N$4735 N$8956 N$8960 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1809 N$8833 N$6974 N$6849 N$6851 "Waveguide Crossing" sch_x=124 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1810 N$6976 N$6978 N$6853 N$6855 "Waveguide Crossing" sch_x=124 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1811 N$6980 N$6982 N$6857 N$6859 "Waveguide Crossing" sch_x=124 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1812 N$6984 N$6986 N$6861 N$6863 "Waveguide Crossing" sch_x=124 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1813 N$6988 N$6990 N$6865 N$6867 "Waveguide Crossing" sch_x=124 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1814 N$6992 N$6994 N$6869 N$6871 "Waveguide Crossing" sch_x=124 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1815 N$6996 N$6998 N$6873 N$6875 "Waveguide Crossing" sch_x=124 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1816 N$7000 N$7002 N$6877 N$6879 "Waveguide Crossing" sch_x=124 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1817 N$7004 N$7006 N$6881 N$6883 "Waveguide Crossing" sch_x=124 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1818 N$7008 N$7010 N$6885 N$6887 "Waveguide Crossing" sch_x=124 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1819 N$7012 N$7014 N$6889 N$6891 "Waveguide Crossing" sch_x=124 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1820 N$7016 N$7018 N$6893 N$6895 "Waveguide Crossing" sch_x=124 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1821 N$7020 N$7022 N$6897 N$6899 "Waveguide Crossing" sch_x=124 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1822 N$7024 N$7026 N$6901 N$6903 "Waveguide Crossing" sch_x=124 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1823 N$7028 N$7030 N$6905 N$6907 "Waveguide Crossing" sch_x=124 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1824 N$7032 N$7034 N$6909 N$6911 "Waveguide Crossing" sch_x=124 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1825 N$7036 N$7038 N$6913 N$6915 "Waveguide Crossing" sch_x=124 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1826 N$7040 N$7042 N$6917 N$6919 "Waveguide Crossing" sch_x=124 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1827 N$7044 N$7046 N$6921 N$6923 "Waveguide Crossing" sch_x=124 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1828 N$7048 N$7050 N$6925 N$6927 "Waveguide Crossing" sch_x=124 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1829 N$7052 N$7054 N$6929 N$6931 "Waveguide Crossing" sch_x=124 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1830 N$7056 N$7058 N$6933 N$6935 "Waveguide Crossing" sch_x=124 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1831 N$7060 N$7062 N$6937 N$6939 "Waveguide Crossing" sch_x=124 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1832 N$7064 N$7066 N$6941 N$6943 "Waveguide Crossing" sch_x=124 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1833 N$7068 N$7070 N$6945 N$6947 "Waveguide Crossing" sch_x=124 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1834 N$7072 N$7074 N$6949 N$6951 "Waveguide Crossing" sch_x=124 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1835 N$7076 N$7078 N$6953 N$6955 "Waveguide Crossing" sch_x=124 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1836 N$7080 N$7082 N$6957 N$6959 "Waveguide Crossing" sch_x=124 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1837 N$7084 N$7086 N$6961 N$6963 "Waveguide Crossing" sch_x=124 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1838 N$7088 N$7090 N$6965 N$6967 "Waveguide Crossing" sch_x=124 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1839 N$7092 N$8955 N$6969 N$6971 "Waveguide Crossing" sch_x=124 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1840 N$8835 N$7094 N$6973 N$6975 "Waveguide Crossing" sch_x=122 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1841 N$7096 N$7098 N$6977 N$6979 "Waveguide Crossing" sch_x=122 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1842 N$7100 N$7102 N$6981 N$6983 "Waveguide Crossing" sch_x=122 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1843 N$7104 N$7106 N$6985 N$6987 "Waveguide Crossing" sch_x=122 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1844 N$7108 N$7110 N$6989 N$6991 "Waveguide Crossing" sch_x=122 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1845 N$7112 N$7114 N$6993 N$6995 "Waveguide Crossing" sch_x=122 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1846 N$7116 N$7118 N$6997 N$6999 "Waveguide Crossing" sch_x=122 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1847 N$7120 N$7122 N$7001 N$7003 "Waveguide Crossing" sch_x=122 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1848 N$7124 N$7126 N$7005 N$7007 "Waveguide Crossing" sch_x=122 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1849 N$7128 N$7130 N$7009 N$7011 "Waveguide Crossing" sch_x=122 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1850 N$7132 N$7134 N$7013 N$7015 "Waveguide Crossing" sch_x=122 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1851 N$7136 N$7138 N$7017 N$7019 "Waveguide Crossing" sch_x=122 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1852 N$7140 N$7142 N$7021 N$7023 "Waveguide Crossing" sch_x=122 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1853 N$7144 N$7146 N$7025 N$7027 "Waveguide Crossing" sch_x=122 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1854 N$7148 N$7150 N$7029 N$7031 "Waveguide Crossing" sch_x=122 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1855 N$7152 N$7154 N$7033 N$7035 "Waveguide Crossing" sch_x=122 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1856 N$7156 N$7158 N$7037 N$7039 "Waveguide Crossing" sch_x=122 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1857 N$7160 N$7162 N$7041 N$7043 "Waveguide Crossing" sch_x=122 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1858 N$7164 N$7166 N$7045 N$7047 "Waveguide Crossing" sch_x=122 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1859 N$7168 N$7170 N$7049 N$7051 "Waveguide Crossing" sch_x=122 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1860 N$7172 N$7174 N$7053 N$7055 "Waveguide Crossing" sch_x=122 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1861 N$7176 N$7178 N$7057 N$7059 "Waveguide Crossing" sch_x=122 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1862 N$7180 N$7182 N$7061 N$7063 "Waveguide Crossing" sch_x=122 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1863 N$7184 N$7186 N$7065 N$7067 "Waveguide Crossing" sch_x=122 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1864 N$7188 N$7190 N$7069 N$7071 "Waveguide Crossing" sch_x=122 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1865 N$7192 N$7194 N$7073 N$7075 "Waveguide Crossing" sch_x=122 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1866 N$7196 N$7198 N$7077 N$7079 "Waveguide Crossing" sch_x=122 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1867 N$7200 N$7202 N$7081 N$7083 "Waveguide Crossing" sch_x=122 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1868 N$7204 N$7206 N$7085 N$7087 "Waveguide Crossing" sch_x=122 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1869 N$7208 N$8953 N$7089 N$7091 "Waveguide Crossing" sch_x=122 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1870 N$8837 N$7210 N$7093 N$7095 "Waveguide Crossing" sch_x=120 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1871 N$7212 N$7214 N$7097 N$7099 "Waveguide Crossing" sch_x=120 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1872 N$7216 N$7218 N$7101 N$7103 "Waveguide Crossing" sch_x=120 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1873 N$7220 N$7222 N$7105 N$7107 "Waveguide Crossing" sch_x=120 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1874 N$7224 N$7226 N$7109 N$7111 "Waveguide Crossing" sch_x=120 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1875 N$7228 N$7230 N$7113 N$7115 "Waveguide Crossing" sch_x=120 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1876 N$7232 N$7234 N$7117 N$7119 "Waveguide Crossing" sch_x=120 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1877 N$7236 N$7238 N$7121 N$7123 "Waveguide Crossing" sch_x=120 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1878 N$7240 N$7242 N$7125 N$7127 "Waveguide Crossing" sch_x=120 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1879 N$7244 N$7246 N$7129 N$7131 "Waveguide Crossing" sch_x=120 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1880 N$7248 N$7250 N$7133 N$7135 "Waveguide Crossing" sch_x=120 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1881 N$7252 N$7254 N$7137 N$7139 "Waveguide Crossing" sch_x=120 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1882 N$7256 N$7258 N$7141 N$7143 "Waveguide Crossing" sch_x=120 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1883 N$7260 N$7262 N$7145 N$7147 "Waveguide Crossing" sch_x=120 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1884 N$7264 N$7266 N$7149 N$7151 "Waveguide Crossing" sch_x=120 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1885 N$7268 N$7270 N$7153 N$7155 "Waveguide Crossing" sch_x=120 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1886 N$7272 N$7274 N$7157 N$7159 "Waveguide Crossing" sch_x=120 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1887 N$7276 N$7278 N$7161 N$7163 "Waveguide Crossing" sch_x=120 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1888 N$7280 N$7282 N$7165 N$7167 "Waveguide Crossing" sch_x=120 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1889 N$7284 N$7286 N$7169 N$7171 "Waveguide Crossing" sch_x=120 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1890 N$7288 N$7290 N$7173 N$7175 "Waveguide Crossing" sch_x=120 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1891 N$7292 N$7294 N$7177 N$7179 "Waveguide Crossing" sch_x=120 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1892 N$7296 N$7298 N$7181 N$7183 "Waveguide Crossing" sch_x=120 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1893 N$7300 N$7302 N$7185 N$7187 "Waveguide Crossing" sch_x=120 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1894 N$7304 N$7306 N$7189 N$7191 "Waveguide Crossing" sch_x=120 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1895 N$7308 N$7310 N$7193 N$7195 "Waveguide Crossing" sch_x=120 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1896 N$7312 N$7314 N$7197 N$7199 "Waveguide Crossing" sch_x=120 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1897 N$7316 N$7318 N$7201 N$7203 "Waveguide Crossing" sch_x=120 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1898 N$7320 N$8951 N$7205 N$7207 "Waveguide Crossing" sch_x=120 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1899 N$8839 N$7322 N$7209 N$7211 "Waveguide Crossing" sch_x=118 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1900 N$7324 N$7326 N$7213 N$7215 "Waveguide Crossing" sch_x=118 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1901 N$7328 N$7330 N$7217 N$7219 "Waveguide Crossing" sch_x=118 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1902 N$7332 N$7334 N$7221 N$7223 "Waveguide Crossing" sch_x=118 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1903 N$7336 N$7338 N$7225 N$7227 "Waveguide Crossing" sch_x=118 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1904 N$7340 N$7342 N$7229 N$7231 "Waveguide Crossing" sch_x=118 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1905 N$7344 N$7346 N$7233 N$7235 "Waveguide Crossing" sch_x=118 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1906 N$7348 N$7350 N$7237 N$7239 "Waveguide Crossing" sch_x=118 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1907 N$7352 N$7354 N$7241 N$7243 "Waveguide Crossing" sch_x=118 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1908 N$7356 N$7358 N$7245 N$7247 "Waveguide Crossing" sch_x=118 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1909 N$7360 N$7362 N$7249 N$7251 "Waveguide Crossing" sch_x=118 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1910 N$7364 N$7366 N$7253 N$7255 "Waveguide Crossing" sch_x=118 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1911 N$7368 N$7370 N$7257 N$7259 "Waveguide Crossing" sch_x=118 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1912 N$7372 N$7374 N$7261 N$7263 "Waveguide Crossing" sch_x=118 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1913 N$7376 N$7378 N$7265 N$7267 "Waveguide Crossing" sch_x=118 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1914 N$7380 N$7382 N$7269 N$7271 "Waveguide Crossing" sch_x=118 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1915 N$7384 N$7386 N$7273 N$7275 "Waveguide Crossing" sch_x=118 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1916 N$7388 N$7390 N$7277 N$7279 "Waveguide Crossing" sch_x=118 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1917 N$7392 N$7394 N$7281 N$7283 "Waveguide Crossing" sch_x=118 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1918 N$7396 N$7398 N$7285 N$7287 "Waveguide Crossing" sch_x=118 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1919 N$7400 N$7402 N$7289 N$7291 "Waveguide Crossing" sch_x=118 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1920 N$7404 N$7406 N$7293 N$7295 "Waveguide Crossing" sch_x=118 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1921 N$7408 N$7410 N$7297 N$7299 "Waveguide Crossing" sch_x=118 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1922 N$7412 N$7414 N$7301 N$7303 "Waveguide Crossing" sch_x=118 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1923 N$7416 N$7418 N$7305 N$7307 "Waveguide Crossing" sch_x=118 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1924 N$7420 N$7422 N$7309 N$7311 "Waveguide Crossing" sch_x=118 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1925 N$7424 N$7426 N$7313 N$7315 "Waveguide Crossing" sch_x=118 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1926 N$7428 N$8949 N$7317 N$7319 "Waveguide Crossing" sch_x=118 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1927 N$8841 N$7430 N$7321 N$7323 "Waveguide Crossing" sch_x=116 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1928 N$7432 N$7434 N$7325 N$7327 "Waveguide Crossing" sch_x=116 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1929 N$7436 N$7438 N$7329 N$7331 "Waveguide Crossing" sch_x=116 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1930 N$7440 N$7442 N$7333 N$7335 "Waveguide Crossing" sch_x=116 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1931 N$7444 N$7446 N$7337 N$7339 "Waveguide Crossing" sch_x=116 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1932 N$7448 N$7450 N$7341 N$7343 "Waveguide Crossing" sch_x=116 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1933 N$7452 N$7454 N$7345 N$7347 "Waveguide Crossing" sch_x=116 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1934 N$7456 N$7458 N$7349 N$7351 "Waveguide Crossing" sch_x=116 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1935 N$7460 N$7462 N$7353 N$7355 "Waveguide Crossing" sch_x=116 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1936 N$7464 N$7466 N$7357 N$7359 "Waveguide Crossing" sch_x=116 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1937 N$7468 N$7470 N$7361 N$7363 "Waveguide Crossing" sch_x=116 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1938 N$7472 N$7474 N$7365 N$7367 "Waveguide Crossing" sch_x=116 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1939 N$7476 N$7478 N$7369 N$7371 "Waveguide Crossing" sch_x=116 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1940 N$7480 N$7482 N$7373 N$7375 "Waveguide Crossing" sch_x=116 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1941 N$7484 N$7486 N$7377 N$7379 "Waveguide Crossing" sch_x=116 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1942 N$7488 N$7490 N$7381 N$7383 "Waveguide Crossing" sch_x=116 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1943 N$7492 N$7494 N$7385 N$7387 "Waveguide Crossing" sch_x=116 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1944 N$7496 N$7498 N$7389 N$7391 "Waveguide Crossing" sch_x=116 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1945 N$7500 N$7502 N$7393 N$7395 "Waveguide Crossing" sch_x=116 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1946 N$7504 N$7506 N$7397 N$7399 "Waveguide Crossing" sch_x=116 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1947 N$7508 N$7510 N$7401 N$7403 "Waveguide Crossing" sch_x=116 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1948 N$7512 N$7514 N$7405 N$7407 "Waveguide Crossing" sch_x=116 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1949 N$7516 N$7518 N$7409 N$7411 "Waveguide Crossing" sch_x=116 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1950 N$7520 N$7522 N$7413 N$7415 "Waveguide Crossing" sch_x=116 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1951 N$7524 N$7526 N$7417 N$7419 "Waveguide Crossing" sch_x=116 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1952 N$7528 N$7530 N$7421 N$7423 "Waveguide Crossing" sch_x=116 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1953 N$7532 N$8947 N$7425 N$7427 "Waveguide Crossing" sch_x=116 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1954 N$8843 N$7534 N$7429 N$7431 "Waveguide Crossing" sch_x=114 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1955 N$7536 N$7538 N$7433 N$7435 "Waveguide Crossing" sch_x=114 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1956 N$7540 N$7542 N$7437 N$7439 "Waveguide Crossing" sch_x=114 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1957 N$7544 N$7546 N$7441 N$7443 "Waveguide Crossing" sch_x=114 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1958 N$7548 N$7550 N$7445 N$7447 "Waveguide Crossing" sch_x=114 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1959 N$7552 N$7554 N$7449 N$7451 "Waveguide Crossing" sch_x=114 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1960 N$7556 N$7558 N$7453 N$7455 "Waveguide Crossing" sch_x=114 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1961 N$7560 N$7562 N$7457 N$7459 "Waveguide Crossing" sch_x=114 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1962 N$7564 N$7566 N$7461 N$7463 "Waveguide Crossing" sch_x=114 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1963 N$7568 N$7570 N$7465 N$7467 "Waveguide Crossing" sch_x=114 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1964 N$7572 N$7574 N$7469 N$7471 "Waveguide Crossing" sch_x=114 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1965 N$7576 N$7578 N$7473 N$7475 "Waveguide Crossing" sch_x=114 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1966 N$7580 N$7582 N$7477 N$7479 "Waveguide Crossing" sch_x=114 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1967 N$7584 N$7586 N$7481 N$7483 "Waveguide Crossing" sch_x=114 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1968 N$7588 N$7590 N$7485 N$7487 "Waveguide Crossing" sch_x=114 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1969 N$7592 N$7594 N$7489 N$7491 "Waveguide Crossing" sch_x=114 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1970 N$7596 N$7598 N$7493 N$7495 "Waveguide Crossing" sch_x=114 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1971 N$7600 N$7602 N$7497 N$7499 "Waveguide Crossing" sch_x=114 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1972 N$7604 N$7606 N$7501 N$7503 "Waveguide Crossing" sch_x=114 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1973 N$7608 N$7610 N$7505 N$7507 "Waveguide Crossing" sch_x=114 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1974 N$7612 N$7614 N$7509 N$7511 "Waveguide Crossing" sch_x=114 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1975 N$7616 N$7618 N$7513 N$7515 "Waveguide Crossing" sch_x=114 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1976 N$7620 N$7622 N$7517 N$7519 "Waveguide Crossing" sch_x=114 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1977 N$7624 N$7626 N$7521 N$7523 "Waveguide Crossing" sch_x=114 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1978 N$7628 N$7630 N$7525 N$7527 "Waveguide Crossing" sch_x=114 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1979 N$7632 N$8945 N$7529 N$7531 "Waveguide Crossing" sch_x=114 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1980 N$8845 N$7634 N$7533 N$7535 "Waveguide Crossing" sch_x=112 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1981 N$7636 N$7638 N$7537 N$7539 "Waveguide Crossing" sch_x=112 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1982 N$7640 N$7642 N$7541 N$7543 "Waveguide Crossing" sch_x=112 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1983 N$7644 N$7646 N$7545 N$7547 "Waveguide Crossing" sch_x=112 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1984 N$7648 N$7650 N$7549 N$7551 "Waveguide Crossing" sch_x=112 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1985 N$7652 N$7654 N$7553 N$7555 "Waveguide Crossing" sch_x=112 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1986 N$7656 N$7658 N$7557 N$7559 "Waveguide Crossing" sch_x=112 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1987 N$7660 N$7662 N$7561 N$7563 "Waveguide Crossing" sch_x=112 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1988 N$7664 N$7666 N$7565 N$7567 "Waveguide Crossing" sch_x=112 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1989 N$7668 N$7670 N$7569 N$7571 "Waveguide Crossing" sch_x=112 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1990 N$7672 N$7674 N$7573 N$7575 "Waveguide Crossing" sch_x=112 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1991 N$7676 N$7678 N$7577 N$7579 "Waveguide Crossing" sch_x=112 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1992 N$7680 N$7682 N$7581 N$7583 "Waveguide Crossing" sch_x=112 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1993 N$7684 N$7686 N$7585 N$7587 "Waveguide Crossing" sch_x=112 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1994 N$7688 N$7690 N$7589 N$7591 "Waveguide Crossing" sch_x=112 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1995 N$7692 N$7694 N$7593 N$7595 "Waveguide Crossing" sch_x=112 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1996 N$7696 N$7698 N$7597 N$7599 "Waveguide Crossing" sch_x=112 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1997 N$7700 N$7702 N$7601 N$7603 "Waveguide Crossing" sch_x=112 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1998 N$7704 N$7706 N$7605 N$7607 "Waveguide Crossing" sch_x=112 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1999 N$7708 N$7710 N$7609 N$7611 "Waveguide Crossing" sch_x=112 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2000 N$7712 N$7714 N$7613 N$7615 "Waveguide Crossing" sch_x=112 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2001 N$7716 N$7718 N$7617 N$7619 "Waveguide Crossing" sch_x=112 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2002 N$7720 N$7722 N$7621 N$7623 "Waveguide Crossing" sch_x=112 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2003 N$7724 N$7726 N$7625 N$7627 "Waveguide Crossing" sch_x=112 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2004 N$7728 N$8943 N$7629 N$7631 "Waveguide Crossing" sch_x=112 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2005 N$8847 N$7730 N$7633 N$7635 "Waveguide Crossing" sch_x=110 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2006 N$7732 N$7734 N$7637 N$7639 "Waveguide Crossing" sch_x=110 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2007 N$7736 N$7738 N$7641 N$7643 "Waveguide Crossing" sch_x=110 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2008 N$7740 N$7742 N$7645 N$7647 "Waveguide Crossing" sch_x=110 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2009 N$7744 N$7746 N$7649 N$7651 "Waveguide Crossing" sch_x=110 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2010 N$7748 N$7750 N$7653 N$7655 "Waveguide Crossing" sch_x=110 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2011 N$7752 N$7754 N$7657 N$7659 "Waveguide Crossing" sch_x=110 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2012 N$7756 N$7758 N$7661 N$7663 "Waveguide Crossing" sch_x=110 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2013 N$7760 N$7762 N$7665 N$7667 "Waveguide Crossing" sch_x=110 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2014 N$7764 N$7766 N$7669 N$7671 "Waveguide Crossing" sch_x=110 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2015 N$7768 N$7770 N$7673 N$7675 "Waveguide Crossing" sch_x=110 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2016 N$7772 N$7774 N$7677 N$7679 "Waveguide Crossing" sch_x=110 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2017 N$7776 N$7778 N$7681 N$7683 "Waveguide Crossing" sch_x=110 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2018 N$7780 N$7782 N$7685 N$7687 "Waveguide Crossing" sch_x=110 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2019 N$7784 N$7786 N$7689 N$7691 "Waveguide Crossing" sch_x=110 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2020 N$7788 N$7790 N$7693 N$7695 "Waveguide Crossing" sch_x=110 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2021 N$7792 N$7794 N$7697 N$7699 "Waveguide Crossing" sch_x=110 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2022 N$7796 N$7798 N$7701 N$7703 "Waveguide Crossing" sch_x=110 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2023 N$7800 N$7802 N$7705 N$7707 "Waveguide Crossing" sch_x=110 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2024 N$7804 N$7806 N$7709 N$7711 "Waveguide Crossing" sch_x=110 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2025 N$7808 N$7810 N$7713 N$7715 "Waveguide Crossing" sch_x=110 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2026 N$7812 N$7814 N$7717 N$7719 "Waveguide Crossing" sch_x=110 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2027 N$7816 N$7818 N$7721 N$7723 "Waveguide Crossing" sch_x=110 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2028 N$7820 N$8941 N$7725 N$7727 "Waveguide Crossing" sch_x=110 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2029 N$8849 N$7822 N$7729 N$7731 "Waveguide Crossing" sch_x=108 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2030 N$7824 N$7826 N$7733 N$7735 "Waveguide Crossing" sch_x=108 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2031 N$7828 N$7830 N$7737 N$7739 "Waveguide Crossing" sch_x=108 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2032 N$7832 N$7834 N$7741 N$7743 "Waveguide Crossing" sch_x=108 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2033 N$7836 N$7838 N$7745 N$7747 "Waveguide Crossing" sch_x=108 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2034 N$7840 N$7842 N$7749 N$7751 "Waveguide Crossing" sch_x=108 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2035 N$7844 N$7846 N$7753 N$7755 "Waveguide Crossing" sch_x=108 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2036 N$7848 N$7850 N$7757 N$7759 "Waveguide Crossing" sch_x=108 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2037 N$7852 N$7854 N$7761 N$7763 "Waveguide Crossing" sch_x=108 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2038 N$7856 N$7858 N$7765 N$7767 "Waveguide Crossing" sch_x=108 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2039 N$7860 N$7862 N$7769 N$7771 "Waveguide Crossing" sch_x=108 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2040 N$7864 N$7866 N$7773 N$7775 "Waveguide Crossing" sch_x=108 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2041 N$7868 N$7870 N$7777 N$7779 "Waveguide Crossing" sch_x=108 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2042 N$7872 N$7874 N$7781 N$7783 "Waveguide Crossing" sch_x=108 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2043 N$7876 N$7878 N$7785 N$7787 "Waveguide Crossing" sch_x=108 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2044 N$7880 N$7882 N$7789 N$7791 "Waveguide Crossing" sch_x=108 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2045 N$7884 N$7886 N$7793 N$7795 "Waveguide Crossing" sch_x=108 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2046 N$7888 N$7890 N$7797 N$7799 "Waveguide Crossing" sch_x=108 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2047 N$7892 N$7894 N$7801 N$7803 "Waveguide Crossing" sch_x=108 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2048 N$7896 N$7898 N$7805 N$7807 "Waveguide Crossing" sch_x=108 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2049 N$7900 N$7902 N$7809 N$7811 "Waveguide Crossing" sch_x=108 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2050 N$7904 N$7906 N$7813 N$7815 "Waveguide Crossing" sch_x=108 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2051 N$7908 N$8939 N$7817 N$7819 "Waveguide Crossing" sch_x=108 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2052 N$8851 N$7910 N$7821 N$7823 "Waveguide Crossing" sch_x=106 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2053 N$7912 N$7914 N$7825 N$7827 "Waveguide Crossing" sch_x=106 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2054 N$7916 N$7918 N$7829 N$7831 "Waveguide Crossing" sch_x=106 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2055 N$7920 N$7922 N$7833 N$7835 "Waveguide Crossing" sch_x=106 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2056 N$7924 N$7926 N$7837 N$7839 "Waveguide Crossing" sch_x=106 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2057 N$7928 N$7930 N$7841 N$7843 "Waveguide Crossing" sch_x=106 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2058 N$7932 N$7934 N$7845 N$7847 "Waveguide Crossing" sch_x=106 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2059 N$7936 N$7938 N$7849 N$7851 "Waveguide Crossing" sch_x=106 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2060 N$7940 N$7942 N$7853 N$7855 "Waveguide Crossing" sch_x=106 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2061 N$7944 N$7946 N$7857 N$7859 "Waveguide Crossing" sch_x=106 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2062 N$7948 N$7950 N$7861 N$7863 "Waveguide Crossing" sch_x=106 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2063 N$7952 N$7954 N$7865 N$7867 "Waveguide Crossing" sch_x=106 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2064 N$7956 N$7958 N$7869 N$7871 "Waveguide Crossing" sch_x=106 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2065 N$7960 N$7962 N$7873 N$7875 "Waveguide Crossing" sch_x=106 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2066 N$7964 N$7966 N$7877 N$7879 "Waveguide Crossing" sch_x=106 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2067 N$7968 N$7970 N$7881 N$7883 "Waveguide Crossing" sch_x=106 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2068 N$7972 N$7974 N$7885 N$7887 "Waveguide Crossing" sch_x=106 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2069 N$7976 N$7978 N$7889 N$7891 "Waveguide Crossing" sch_x=106 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2070 N$7980 N$7982 N$7893 N$7895 "Waveguide Crossing" sch_x=106 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2071 N$7984 N$7986 N$7897 N$7899 "Waveguide Crossing" sch_x=106 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2072 N$7988 N$7990 N$7901 N$7903 "Waveguide Crossing" sch_x=106 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2073 N$7992 N$8937 N$7905 N$7907 "Waveguide Crossing" sch_x=106 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2074 N$8853 N$7994 N$7909 N$7911 "Waveguide Crossing" sch_x=104 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2075 N$7996 N$7998 N$7913 N$7915 "Waveguide Crossing" sch_x=104 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2076 N$8000 N$8002 N$7917 N$7919 "Waveguide Crossing" sch_x=104 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2077 N$8004 N$8006 N$7921 N$7923 "Waveguide Crossing" sch_x=104 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2078 N$8008 N$8010 N$7925 N$7927 "Waveguide Crossing" sch_x=104 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2079 N$8012 N$8014 N$7929 N$7931 "Waveguide Crossing" sch_x=104 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2080 N$8016 N$8018 N$7933 N$7935 "Waveguide Crossing" sch_x=104 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2081 N$8020 N$8022 N$7937 N$7939 "Waveguide Crossing" sch_x=104 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2082 N$8024 N$8026 N$7941 N$7943 "Waveguide Crossing" sch_x=104 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2083 N$8028 N$8030 N$7945 N$7947 "Waveguide Crossing" sch_x=104 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2084 N$8032 N$8034 N$7949 N$7951 "Waveguide Crossing" sch_x=104 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2085 N$8036 N$8038 N$7953 N$7955 "Waveguide Crossing" sch_x=104 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2086 N$8040 N$8042 N$7957 N$7959 "Waveguide Crossing" sch_x=104 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2087 N$8044 N$8046 N$7961 N$7963 "Waveguide Crossing" sch_x=104 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2088 N$8048 N$8050 N$7965 N$7967 "Waveguide Crossing" sch_x=104 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2089 N$8052 N$8054 N$7969 N$7971 "Waveguide Crossing" sch_x=104 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2090 N$8056 N$8058 N$7973 N$7975 "Waveguide Crossing" sch_x=104 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2091 N$8060 N$8062 N$7977 N$7979 "Waveguide Crossing" sch_x=104 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2092 N$8064 N$8066 N$7981 N$7983 "Waveguide Crossing" sch_x=104 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2093 N$8068 N$8070 N$7985 N$7987 "Waveguide Crossing" sch_x=104 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2094 N$8072 N$8935 N$7989 N$7991 "Waveguide Crossing" sch_x=104 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2095 N$8855 N$8074 N$7993 N$7995 "Waveguide Crossing" sch_x=102 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2096 N$8076 N$8078 N$7997 N$7999 "Waveguide Crossing" sch_x=102 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2097 N$8080 N$8082 N$8001 N$8003 "Waveguide Crossing" sch_x=102 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2098 N$8084 N$8086 N$8005 N$8007 "Waveguide Crossing" sch_x=102 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2099 N$8088 N$8090 N$8009 N$8011 "Waveguide Crossing" sch_x=102 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2100 N$8092 N$8094 N$8013 N$8015 "Waveguide Crossing" sch_x=102 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2101 N$8096 N$8098 N$8017 N$8019 "Waveguide Crossing" sch_x=102 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2102 N$8100 N$8102 N$8021 N$8023 "Waveguide Crossing" sch_x=102 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2103 N$8104 N$8106 N$8025 N$8027 "Waveguide Crossing" sch_x=102 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2104 N$8108 N$8110 N$8029 N$8031 "Waveguide Crossing" sch_x=102 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2105 N$8112 N$8114 N$8033 N$8035 "Waveguide Crossing" sch_x=102 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2106 N$8116 N$8118 N$8037 N$8039 "Waveguide Crossing" sch_x=102 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2107 N$8120 N$8122 N$8041 N$8043 "Waveguide Crossing" sch_x=102 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2108 N$8124 N$8126 N$8045 N$8047 "Waveguide Crossing" sch_x=102 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2109 N$8128 N$8130 N$8049 N$8051 "Waveguide Crossing" sch_x=102 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2110 N$8132 N$8134 N$8053 N$8055 "Waveguide Crossing" sch_x=102 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2111 N$8136 N$8138 N$8057 N$8059 "Waveguide Crossing" sch_x=102 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2112 N$8140 N$8142 N$8061 N$8063 "Waveguide Crossing" sch_x=102 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2113 N$8144 N$8146 N$8065 N$8067 "Waveguide Crossing" sch_x=102 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2114 N$8148 N$8933 N$8069 N$8071 "Waveguide Crossing" sch_x=102 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2115 N$8857 N$8150 N$8073 N$8075 "Waveguide Crossing" sch_x=100 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2116 N$8152 N$8154 N$8077 N$8079 "Waveguide Crossing" sch_x=100 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2117 N$8156 N$8158 N$8081 N$8083 "Waveguide Crossing" sch_x=100 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2118 N$8160 N$8162 N$8085 N$8087 "Waveguide Crossing" sch_x=100 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2119 N$8164 N$8166 N$8089 N$8091 "Waveguide Crossing" sch_x=100 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2120 N$8168 N$8170 N$8093 N$8095 "Waveguide Crossing" sch_x=100 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2121 N$8172 N$8174 N$8097 N$8099 "Waveguide Crossing" sch_x=100 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2122 N$8176 N$8178 N$8101 N$8103 "Waveguide Crossing" sch_x=100 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2123 N$8180 N$8182 N$8105 N$8107 "Waveguide Crossing" sch_x=100 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2124 N$8184 N$8186 N$8109 N$8111 "Waveguide Crossing" sch_x=100 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2125 N$8188 N$8190 N$8113 N$8115 "Waveguide Crossing" sch_x=100 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2126 N$8192 N$8194 N$8117 N$8119 "Waveguide Crossing" sch_x=100 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2127 N$8196 N$8198 N$8121 N$8123 "Waveguide Crossing" sch_x=100 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2128 N$8200 N$8202 N$8125 N$8127 "Waveguide Crossing" sch_x=100 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2129 N$8204 N$8206 N$8129 N$8131 "Waveguide Crossing" sch_x=100 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2130 N$8208 N$8210 N$8133 N$8135 "Waveguide Crossing" sch_x=100 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2131 N$8212 N$8214 N$8137 N$8139 "Waveguide Crossing" sch_x=100 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2132 N$8216 N$8218 N$8141 N$8143 "Waveguide Crossing" sch_x=100 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2133 N$8220 N$8931 N$8145 N$8147 "Waveguide Crossing" sch_x=100 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2134 N$8859 N$8222 N$8149 N$8151 "Waveguide Crossing" sch_x=98 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2135 N$8224 N$8226 N$8153 N$8155 "Waveguide Crossing" sch_x=98 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2136 N$8228 N$8230 N$8157 N$8159 "Waveguide Crossing" sch_x=98 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2137 N$8232 N$8234 N$8161 N$8163 "Waveguide Crossing" sch_x=98 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2138 N$8236 N$8238 N$8165 N$8167 "Waveguide Crossing" sch_x=98 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2139 N$8240 N$8242 N$8169 N$8171 "Waveguide Crossing" sch_x=98 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2140 N$8244 N$8246 N$8173 N$8175 "Waveguide Crossing" sch_x=98 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2141 N$8248 N$8250 N$8177 N$8179 "Waveguide Crossing" sch_x=98 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2142 N$8252 N$8254 N$8181 N$8183 "Waveguide Crossing" sch_x=98 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2143 N$8256 N$8258 N$8185 N$8187 "Waveguide Crossing" sch_x=98 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2144 N$8260 N$8262 N$8189 N$8191 "Waveguide Crossing" sch_x=98 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2145 N$8264 N$8266 N$8193 N$8195 "Waveguide Crossing" sch_x=98 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2146 N$8268 N$8270 N$8197 N$8199 "Waveguide Crossing" sch_x=98 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2147 N$8272 N$8274 N$8201 N$8203 "Waveguide Crossing" sch_x=98 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2148 N$8276 N$8278 N$8205 N$8207 "Waveguide Crossing" sch_x=98 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2149 N$8280 N$8282 N$8209 N$8211 "Waveguide Crossing" sch_x=98 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2150 N$8284 N$8286 N$8213 N$8215 "Waveguide Crossing" sch_x=98 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2151 N$8288 N$8929 N$8217 N$8219 "Waveguide Crossing" sch_x=98 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2152 N$8861 N$8290 N$8221 N$8223 "Waveguide Crossing" sch_x=96 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2153 N$8292 N$8294 N$8225 N$8227 "Waveguide Crossing" sch_x=96 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2154 N$8296 N$8298 N$8229 N$8231 "Waveguide Crossing" sch_x=96 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2155 N$8300 N$8302 N$8233 N$8235 "Waveguide Crossing" sch_x=96 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2156 N$8304 N$8306 N$8237 N$8239 "Waveguide Crossing" sch_x=96 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2157 N$8308 N$8310 N$8241 N$8243 "Waveguide Crossing" sch_x=96 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2158 N$8312 N$8314 N$8245 N$8247 "Waveguide Crossing" sch_x=96 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2159 N$8316 N$8318 N$8249 N$8251 "Waveguide Crossing" sch_x=96 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2160 N$8320 N$8322 N$8253 N$8255 "Waveguide Crossing" sch_x=96 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2161 N$8324 N$8326 N$8257 N$8259 "Waveguide Crossing" sch_x=96 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2162 N$8328 N$8330 N$8261 N$8263 "Waveguide Crossing" sch_x=96 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2163 N$8332 N$8334 N$8265 N$8267 "Waveguide Crossing" sch_x=96 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2164 N$8336 N$8338 N$8269 N$8271 "Waveguide Crossing" sch_x=96 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2165 N$8340 N$8342 N$8273 N$8275 "Waveguide Crossing" sch_x=96 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2166 N$8344 N$8346 N$8277 N$8279 "Waveguide Crossing" sch_x=96 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2167 N$8348 N$8350 N$8281 N$8283 "Waveguide Crossing" sch_x=96 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2168 N$8352 N$8927 N$8285 N$8287 "Waveguide Crossing" sch_x=96 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2169 N$8863 N$8354 N$8289 N$8291 "Waveguide Crossing" sch_x=94 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2170 N$8356 N$8358 N$8293 N$8295 "Waveguide Crossing" sch_x=94 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2171 N$8360 N$8362 N$8297 N$8299 "Waveguide Crossing" sch_x=94 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2172 N$8364 N$8366 N$8301 N$8303 "Waveguide Crossing" sch_x=94 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2173 N$8368 N$8370 N$8305 N$8307 "Waveguide Crossing" sch_x=94 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2174 N$8372 N$8374 N$8309 N$8311 "Waveguide Crossing" sch_x=94 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2175 N$8376 N$8378 N$8313 N$8315 "Waveguide Crossing" sch_x=94 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2176 N$8380 N$8382 N$8317 N$8319 "Waveguide Crossing" sch_x=94 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2177 N$8384 N$8386 N$8321 N$8323 "Waveguide Crossing" sch_x=94 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2178 N$8388 N$8390 N$8325 N$8327 "Waveguide Crossing" sch_x=94 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2179 N$8392 N$8394 N$8329 N$8331 "Waveguide Crossing" sch_x=94 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2180 N$8396 N$8398 N$8333 N$8335 "Waveguide Crossing" sch_x=94 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2181 N$8400 N$8402 N$8337 N$8339 "Waveguide Crossing" sch_x=94 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2182 N$8404 N$8406 N$8341 N$8343 "Waveguide Crossing" sch_x=94 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2183 N$8408 N$8410 N$8345 N$8347 "Waveguide Crossing" sch_x=94 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2184 N$8412 N$8925 N$8349 N$8351 "Waveguide Crossing" sch_x=94 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2185 N$8865 N$8414 N$8353 N$8355 "Waveguide Crossing" sch_x=92 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2186 N$8416 N$8418 N$8357 N$8359 "Waveguide Crossing" sch_x=92 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2187 N$8420 N$8422 N$8361 N$8363 "Waveguide Crossing" sch_x=92 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2188 N$8424 N$8426 N$8365 N$8367 "Waveguide Crossing" sch_x=92 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2189 N$8428 N$8430 N$8369 N$8371 "Waveguide Crossing" sch_x=92 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2190 N$8432 N$8434 N$8373 N$8375 "Waveguide Crossing" sch_x=92 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2191 N$8436 N$8438 N$8377 N$8379 "Waveguide Crossing" sch_x=92 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2192 N$8440 N$8442 N$8381 N$8383 "Waveguide Crossing" sch_x=92 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2193 N$8444 N$8446 N$8385 N$8387 "Waveguide Crossing" sch_x=92 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2194 N$8448 N$8450 N$8389 N$8391 "Waveguide Crossing" sch_x=92 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2195 N$8452 N$8454 N$8393 N$8395 "Waveguide Crossing" sch_x=92 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2196 N$8456 N$8458 N$8397 N$8399 "Waveguide Crossing" sch_x=92 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2197 N$8460 N$8462 N$8401 N$8403 "Waveguide Crossing" sch_x=92 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2198 N$8464 N$8466 N$8405 N$8407 "Waveguide Crossing" sch_x=92 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2199 N$8468 N$8923 N$8409 N$8411 "Waveguide Crossing" sch_x=92 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2200 N$8867 N$8470 N$8413 N$8415 "Waveguide Crossing" sch_x=90 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2201 N$8472 N$8474 N$8417 N$8419 "Waveguide Crossing" sch_x=90 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2202 N$8476 N$8478 N$8421 N$8423 "Waveguide Crossing" sch_x=90 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2203 N$8480 N$8482 N$8425 N$8427 "Waveguide Crossing" sch_x=90 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2204 N$8484 N$8486 N$8429 N$8431 "Waveguide Crossing" sch_x=90 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2205 N$8488 N$8490 N$8433 N$8435 "Waveguide Crossing" sch_x=90 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2206 N$8492 N$8494 N$8437 N$8439 "Waveguide Crossing" sch_x=90 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2207 N$8496 N$8498 N$8441 N$8443 "Waveguide Crossing" sch_x=90 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2208 N$8500 N$8502 N$8445 N$8447 "Waveguide Crossing" sch_x=90 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2209 N$8504 N$8506 N$8449 N$8451 "Waveguide Crossing" sch_x=90 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2210 N$8508 N$8510 N$8453 N$8455 "Waveguide Crossing" sch_x=90 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2211 N$8512 N$8514 N$8457 N$8459 "Waveguide Crossing" sch_x=90 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2212 N$8516 N$8518 N$8461 N$8463 "Waveguide Crossing" sch_x=90 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2213 N$8520 N$8921 N$8465 N$8467 "Waveguide Crossing" sch_x=90 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2214 N$8869 N$8522 N$8469 N$8471 "Waveguide Crossing" sch_x=88 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2215 N$8524 N$8526 N$8473 N$8475 "Waveguide Crossing" sch_x=88 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2216 N$8528 N$8530 N$8477 N$8479 "Waveguide Crossing" sch_x=88 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2217 N$8532 N$8534 N$8481 N$8483 "Waveguide Crossing" sch_x=88 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2218 N$8536 N$8538 N$8485 N$8487 "Waveguide Crossing" sch_x=88 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2219 N$8540 N$8542 N$8489 N$8491 "Waveguide Crossing" sch_x=88 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2220 N$8544 N$8546 N$8493 N$8495 "Waveguide Crossing" sch_x=88 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2221 N$8548 N$8550 N$8497 N$8499 "Waveguide Crossing" sch_x=88 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2222 N$8552 N$8554 N$8501 N$8503 "Waveguide Crossing" sch_x=88 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2223 N$8556 N$8558 N$8505 N$8507 "Waveguide Crossing" sch_x=88 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2224 N$8560 N$8562 N$8509 N$8511 "Waveguide Crossing" sch_x=88 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2225 N$8564 N$8566 N$8513 N$8515 "Waveguide Crossing" sch_x=88 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2226 N$8568 N$8919 N$8517 N$8519 "Waveguide Crossing" sch_x=88 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2227 N$8871 N$8570 N$8521 N$8523 "Waveguide Crossing" sch_x=86 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2228 N$8572 N$8574 N$8525 N$8527 "Waveguide Crossing" sch_x=86 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2229 N$8576 N$8578 N$8529 N$8531 "Waveguide Crossing" sch_x=86 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2230 N$8580 N$8582 N$8533 N$8535 "Waveguide Crossing" sch_x=86 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2231 N$8584 N$8586 N$8537 N$8539 "Waveguide Crossing" sch_x=86 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2232 N$8588 N$8590 N$8541 N$8543 "Waveguide Crossing" sch_x=86 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2233 N$8592 N$8594 N$8545 N$8547 "Waveguide Crossing" sch_x=86 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2234 N$8596 N$8598 N$8549 N$8551 "Waveguide Crossing" sch_x=86 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2235 N$8600 N$8602 N$8553 N$8555 "Waveguide Crossing" sch_x=86 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2236 N$8604 N$8606 N$8557 N$8559 "Waveguide Crossing" sch_x=86 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2237 N$8608 N$8610 N$8561 N$8563 "Waveguide Crossing" sch_x=86 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2238 N$8612 N$8917 N$8565 N$8567 "Waveguide Crossing" sch_x=86 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2239 N$8873 N$8614 N$8569 N$8571 "Waveguide Crossing" sch_x=84 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2240 N$8616 N$8618 N$8573 N$8575 "Waveguide Crossing" sch_x=84 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2241 N$8620 N$8622 N$8577 N$8579 "Waveguide Crossing" sch_x=84 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2242 N$8624 N$8626 N$8581 N$8583 "Waveguide Crossing" sch_x=84 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2243 N$8628 N$8630 N$8585 N$8587 "Waveguide Crossing" sch_x=84 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2244 N$8632 N$8634 N$8589 N$8591 "Waveguide Crossing" sch_x=84 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2245 N$8636 N$8638 N$8593 N$8595 "Waveguide Crossing" sch_x=84 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2246 N$8640 N$8642 N$8597 N$8599 "Waveguide Crossing" sch_x=84 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2247 N$8644 N$8646 N$8601 N$8603 "Waveguide Crossing" sch_x=84 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2248 N$8648 N$8650 N$8605 N$8607 "Waveguide Crossing" sch_x=84 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2249 N$8652 N$8915 N$8609 N$8611 "Waveguide Crossing" sch_x=84 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2250 N$8875 N$8654 N$8613 N$8615 "Waveguide Crossing" sch_x=82 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2251 N$8656 N$8658 N$8617 N$8619 "Waveguide Crossing" sch_x=82 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2252 N$8660 N$8662 N$8621 N$8623 "Waveguide Crossing" sch_x=82 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2253 N$8664 N$8666 N$8625 N$8627 "Waveguide Crossing" sch_x=82 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2254 N$8668 N$8670 N$8629 N$8631 "Waveguide Crossing" sch_x=82 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2255 N$8672 N$8674 N$8633 N$8635 "Waveguide Crossing" sch_x=82 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2256 N$8676 N$8678 N$8637 N$8639 "Waveguide Crossing" sch_x=82 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2257 N$8680 N$8682 N$8641 N$8643 "Waveguide Crossing" sch_x=82 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2258 N$8684 N$8686 N$8645 N$8647 "Waveguide Crossing" sch_x=82 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2259 N$8688 N$8913 N$8649 N$8651 "Waveguide Crossing" sch_x=82 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2260 N$8877 N$8690 N$8653 N$8655 "Waveguide Crossing" sch_x=80 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2261 N$8692 N$8694 N$8657 N$8659 "Waveguide Crossing" sch_x=80 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2262 N$8696 N$8698 N$8661 N$8663 "Waveguide Crossing" sch_x=80 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2263 N$8700 N$8702 N$8665 N$8667 "Waveguide Crossing" sch_x=80 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2264 N$8704 N$8706 N$8669 N$8671 "Waveguide Crossing" sch_x=80 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2265 N$8708 N$8710 N$8673 N$8675 "Waveguide Crossing" sch_x=80 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2266 N$8712 N$8714 N$8677 N$8679 "Waveguide Crossing" sch_x=80 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2267 N$8716 N$8718 N$8681 N$8683 "Waveguide Crossing" sch_x=80 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2268 N$8720 N$8911 N$8685 N$8687 "Waveguide Crossing" sch_x=80 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2269 N$8879 N$8722 N$8689 N$8691 "Waveguide Crossing" sch_x=78 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2270 N$8724 N$8726 N$8693 N$8695 "Waveguide Crossing" sch_x=78 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2271 N$8728 N$8730 N$8697 N$8699 "Waveguide Crossing" sch_x=78 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2272 N$8732 N$8734 N$8701 N$8703 "Waveguide Crossing" sch_x=78 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2273 N$8736 N$8738 N$8705 N$8707 "Waveguide Crossing" sch_x=78 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2274 N$8740 N$8742 N$8709 N$8711 "Waveguide Crossing" sch_x=78 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2275 N$8744 N$8746 N$8713 N$8715 "Waveguide Crossing" sch_x=78 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2276 N$8748 N$8909 N$8717 N$8719 "Waveguide Crossing" sch_x=78 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2277 N$8881 N$8750 N$8721 N$8723 "Waveguide Crossing" sch_x=76 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2278 N$8752 N$8754 N$8725 N$8727 "Waveguide Crossing" sch_x=76 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2279 N$8756 N$8758 N$8729 N$8731 "Waveguide Crossing" sch_x=76 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2280 N$8760 N$8762 N$8733 N$8735 "Waveguide Crossing" sch_x=76 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2281 N$8764 N$8766 N$8737 N$8739 "Waveguide Crossing" sch_x=76 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2282 N$8768 N$8770 N$8741 N$8743 "Waveguide Crossing" sch_x=76 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2283 N$8772 N$8907 N$8745 N$8747 "Waveguide Crossing" sch_x=76 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2284 N$8883 N$8774 N$8749 N$8751 "Waveguide Crossing" sch_x=74 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2285 N$8776 N$8778 N$8753 N$8755 "Waveguide Crossing" sch_x=74 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2286 N$8780 N$8782 N$8757 N$8759 "Waveguide Crossing" sch_x=74 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2287 N$8784 N$8786 N$8761 N$8763 "Waveguide Crossing" sch_x=74 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2288 N$8788 N$8790 N$8765 N$8767 "Waveguide Crossing" sch_x=74 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2289 N$8792 N$8905 N$8769 N$8771 "Waveguide Crossing" sch_x=74 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2290 N$8885 N$8794 N$8773 N$8775 "Waveguide Crossing" sch_x=72 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2291 N$8796 N$8798 N$8777 N$8779 "Waveguide Crossing" sch_x=72 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2292 N$8800 N$8802 N$8781 N$8783 "Waveguide Crossing" sch_x=72 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2293 N$8804 N$8806 N$8785 N$8787 "Waveguide Crossing" sch_x=72 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2294 N$8808 N$8903 N$8789 N$8791 "Waveguide Crossing" sch_x=72 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2295 N$8887 N$8810 N$8793 N$8795 "Waveguide Crossing" sch_x=70 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2296 N$8812 N$8814 N$8797 N$8799 "Waveguide Crossing" sch_x=70 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2297 N$8816 N$8818 N$8801 N$8803 "Waveguide Crossing" sch_x=70 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2298 N$8820 N$8901 N$8805 N$8807 "Waveguide Crossing" sch_x=70 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2299 N$8889 N$8822 N$8809 N$8811 "Waveguide Crossing" sch_x=68 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2300 N$8824 N$8826 N$8813 N$8815 "Waveguide Crossing" sch_x=68 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2301 N$8828 N$8899 N$8817 N$8819 "Waveguide Crossing" sch_x=68 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2302 N$8891 N$8830 N$8821 N$8823 "Waveguide Crossing" sch_x=66 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2303 N$8832 N$8897 N$8825 N$8827 "Waveguide Crossing" sch_x=66 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2304 N$8893 N$8895 N$8829 N$8831 "Waveguide Crossing" sch_x=64 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1777 N$8957 N$6850 N$34558 N$34306 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1778 N$6852 N$6854 N$34308 N$34310 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1779 N$6856 N$6858 N$34312 N$34314 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1780 N$6860 N$6862 N$34316 N$34318 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1781 N$6864 N$6866 N$34320 N$34322 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1782 N$6868 N$6870 N$34324 N$34326 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1783 N$6872 N$6874 N$34328 N$34330 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1784 N$6876 N$6878 N$34332 N$34334 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1785 N$6880 N$6882 N$34336 N$34338 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1786 N$6884 N$6886 N$34340 N$34342 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1787 N$6888 N$6890 N$34344 N$34346 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1788 N$6892 N$6894 N$34348 N$34350 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1789 N$6896 N$6898 N$34352 N$34354 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1790 N$6900 N$6902 N$34356 N$34358 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1791 N$6904 N$6906 N$34360 N$34362 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1792 N$6908 N$6910 N$34364 N$34366 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1793 N$6912 N$6914 N$34368 N$34370 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1794 N$6916 N$6918 N$34372 N$34374 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1795 N$6920 N$6922 N$34376 N$34378 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1796 N$6924 N$6926 N$34380 N$34382 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1797 N$6928 N$6930 N$34384 N$34386 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1798 N$6932 N$6934 N$34388 N$34390 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1799 N$6936 N$6938 N$34392 N$34394 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1800 N$6940 N$6942 N$34396 N$34398 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1801 N$6944 N$6946 N$34400 N$34402 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1802 N$6948 N$6950 N$34404 N$34406 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1803 N$6952 N$6954 N$34408 N$34410 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1804 N$6956 N$6958 N$34412 N$34414 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1805 N$6960 N$6962 N$34416 N$34418 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1806 N$6964 N$6966 N$34420 N$34422 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1807 N$6968 N$6970 N$34424 N$34426 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1808 N$6972 N$8959 N$34428 N$34430 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2305 N$9094 N$9082 N$8961 N$8963 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2306 N$9084 N$9086 N$8965 N$8971 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2307 N$34817 N$8962 N$8973 N$8975 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2308 N$8968 N$34818 N$8977 N$8983 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2309 N$34819 N$8970 N$8985 N$8987 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2310 N$8972 N$34820 N$8989 N$8995 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2311 N$8974 N$8982 N$8997 N$34821 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2312 N$8980 N$8984 N$34822 N$8999 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2313 N$8986 N$8994 N$9001 N$34823 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2314 N$8992 N$8996 N$34824 N$9007 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2315 N$8998 N$9006 N$9134 N$9122 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2316 N$9004 N$9008 N$9124 N$9126 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2317 N$8964 N$8966 N$8967 N$8969 "Waveguide Crossing" sch_x=-4 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2318 N$8976 N$8978 N$8981 N$8979 "Waveguide Crossing" sch_x=0 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2319 N$8988 N$8990 N$8993 N$8991 "Waveguide Crossing" sch_x=0 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2320 N$9000 N$9002 N$9005 N$9003 "Waveguide Crossing" sch_x=4 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2321 N$9088 N$9090 N$9009 N$9011 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2322 N$9092 N$9096 N$9013 N$9019 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2323 N$34825 N$9010 N$9021 N$9023 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2324 N$9016 N$34826 N$9025 N$9031 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2325 N$34827 N$9018 N$9033 N$9035 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2326 N$9020 N$34828 N$9037 N$9043 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2327 N$9022 N$9030 N$9045 N$34829 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2328 N$9028 N$9032 N$34830 N$9047 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2329 N$9034 N$9042 N$9049 N$34831 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2330 N$9040 N$9044 N$34832 N$9055 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2331 N$9046 N$9054 N$9128 N$9130 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2332 N$9052 N$9056 N$9132 N$9136 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2333 N$9012 N$9014 N$9015 N$9017 "Waveguide Crossing" sch_x=-4 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2334 N$9024 N$9026 N$9029 N$9027 "Waveguide Crossing" sch_x=0 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2335 N$9036 N$9038 N$9041 N$9039 "Waveguide Crossing" sch_x=0 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2336 N$9048 N$9050 N$9053 N$9051 "Waveguide Crossing" sch_x=4 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2351 N$9121 N$9110 N$9097 N$9099 "Waveguide Crossing" sch_x=12 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2352 N$9112 N$9114 N$9101 N$9103 "Waveguide Crossing" sch_x=12 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2353 N$9116 N$9131 N$9105 N$9107 "Waveguide Crossing" sch_x=12 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2354 N$9123 N$9118 N$9109 N$9111 "Waveguide Crossing" sch_x=10 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2355 N$9120 N$9129 N$9113 N$9115 "Waveguide Crossing" sch_x=10 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2356 N$9125 N$9127 N$9117 N$9119 "Waveguide Crossing" sch_x=8 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2347 N$9133 N$9098 N$9598 N$9570 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2348 N$9100 N$9102 N$9572 N$9574 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2349 N$9104 N$9106 N$9576 N$9578 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2350 N$9108 N$9135 N$9580 N$9582 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2357 N$9270 N$9258 N$9137 N$9139 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2358 N$9260 N$9262 N$9141 N$9147 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2359 N$34833 N$9138 N$9149 N$9151 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2360 N$9144 N$34834 N$9153 N$9159 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2361 N$34835 N$9146 N$9161 N$9163 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2362 N$9148 N$34836 N$9165 N$9171 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2363 N$9150 N$9158 N$9173 N$34837 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2364 N$9156 N$9160 N$34838 N$9175 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2365 N$9162 N$9170 N$9177 N$34839 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2366 N$9168 N$9172 N$34840 N$9183 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2367 N$9174 N$9182 N$9310 N$9298 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2368 N$9180 N$9184 N$9300 N$9302 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2369 N$9140 N$9142 N$9143 N$9145 "Waveguide Crossing" sch_x=-4 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2370 N$9152 N$9154 N$9157 N$9155 "Waveguide Crossing" sch_x=0 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2371 N$9164 N$9166 N$9169 N$9167 "Waveguide Crossing" sch_x=0 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2372 N$9176 N$9178 N$9181 N$9179 "Waveguide Crossing" sch_x=4 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2373 N$9264 N$9266 N$9185 N$9187 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2374 N$9268 N$9272 N$9189 N$9195 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2375 N$34841 N$9186 N$9197 N$9199 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2376 N$9192 N$34842 N$9201 N$9207 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2377 N$34843 N$9194 N$9209 N$9211 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2378 N$9196 N$34844 N$9213 N$9219 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2379 N$9198 N$9206 N$9221 N$34845 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2380 N$9204 N$9208 N$34846 N$9223 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2381 N$9210 N$9218 N$9225 N$34847 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2382 N$9216 N$9220 N$34848 N$9231 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2383 N$9222 N$9230 N$9304 N$9306 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2384 N$9228 N$9232 N$9308 N$9312 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2385 N$9188 N$9190 N$9191 N$9193 "Waveguide Crossing" sch_x=-4 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2386 N$9200 N$9202 N$9205 N$9203 "Waveguide Crossing" sch_x=0 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2387 N$9212 N$9214 N$9217 N$9215 "Waveguide Crossing" sch_x=0 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2388 N$9224 N$9226 N$9229 N$9227 "Waveguide Crossing" sch_x=4 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2403 N$9297 N$9286 N$9273 N$9275 "Waveguide Crossing" sch_x=12 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2404 N$9288 N$9290 N$9277 N$9279 "Waveguide Crossing" sch_x=12 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2405 N$9292 N$9307 N$9281 N$9283 "Waveguide Crossing" sch_x=12 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2406 N$9299 N$9294 N$9285 N$9287 "Waveguide Crossing" sch_x=10 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2407 N$9296 N$9305 N$9289 N$9291 "Waveguide Crossing" sch_x=10 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2408 N$9301 N$9303 N$9293 N$9295 "Waveguide Crossing" sch_x=8 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2399 N$9309 N$9274 N$9584 N$9586 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2400 N$9276 N$9278 N$9588 N$9590 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2401 N$9280 N$9282 N$9592 N$9594 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2402 N$9284 N$9311 N$9596 N$9600 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2453 N$9569 N$9486 N$9457 N$9459 "Waveguide Crossing" sch_x=28 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2454 N$9488 N$9490 N$9461 N$9463 "Waveguide Crossing" sch_x=28 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2455 N$9492 N$9494 N$9465 N$9467 "Waveguide Crossing" sch_x=28 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2456 N$9496 N$9498 N$9469 N$9471 "Waveguide Crossing" sch_x=28 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2457 N$9500 N$9502 N$9473 N$9475 "Waveguide Crossing" sch_x=28 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2458 N$9504 N$9506 N$9477 N$9479 "Waveguide Crossing" sch_x=28 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2459 N$9508 N$9595 N$9481 N$9483 "Waveguide Crossing" sch_x=28 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2460 N$9571 N$9510 N$9485 N$9487 "Waveguide Crossing" sch_x=26 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2461 N$9512 N$9514 N$9489 N$9491 "Waveguide Crossing" sch_x=26 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2462 N$9516 N$9518 N$9493 N$9495 "Waveguide Crossing" sch_x=26 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2463 N$9520 N$9522 N$9497 N$9499 "Waveguide Crossing" sch_x=26 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2464 N$9524 N$9526 N$9501 N$9503 "Waveguide Crossing" sch_x=26 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2465 N$9528 N$9593 N$9505 N$9507 "Waveguide Crossing" sch_x=26 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2466 N$9573 N$9530 N$9509 N$9511 "Waveguide Crossing" sch_x=24 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2467 N$9532 N$9534 N$9513 N$9515 "Waveguide Crossing" sch_x=24 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2468 N$9536 N$9538 N$9517 N$9519 "Waveguide Crossing" sch_x=24 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2469 N$9540 N$9542 N$9521 N$9523 "Waveguide Crossing" sch_x=24 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2470 N$9544 N$9591 N$9525 N$9527 "Waveguide Crossing" sch_x=24 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2471 N$9575 N$9546 N$9529 N$9531 "Waveguide Crossing" sch_x=22 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2472 N$9548 N$9550 N$9533 N$9535 "Waveguide Crossing" sch_x=22 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2473 N$9552 N$9554 N$9537 N$9539 "Waveguide Crossing" sch_x=22 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2474 N$9556 N$9589 N$9541 N$9543 "Waveguide Crossing" sch_x=22 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2475 N$9577 N$9558 N$9545 N$9547 "Waveguide Crossing" sch_x=20 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2476 N$9560 N$9562 N$9549 N$9551 "Waveguide Crossing" sch_x=20 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2477 N$9564 N$9587 N$9553 N$9555 "Waveguide Crossing" sch_x=20 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2478 N$9579 N$9566 N$9557 N$9559 "Waveguide Crossing" sch_x=18 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2479 N$9568 N$9585 N$9561 N$9563 "Waveguide Crossing" sch_x=18 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2480 N$9581 N$9583 N$9565 N$9567 "Waveguide Crossing" sch_x=16 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2445 N$9597 N$9458 N$11326 N$11266 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2446 N$9460 N$9462 N$11268 N$11270 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2447 N$9464 N$9466 N$11272 N$11274 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2448 N$9468 N$9470 N$11276 N$11278 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2449 N$9472 N$9474 N$11280 N$11282 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2450 N$9476 N$9478 N$11284 N$11286 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2451 N$9480 N$9482 N$11288 N$11290 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2452 N$9484 N$9599 N$11292 N$11294 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2481 N$9734 N$9722 N$9601 N$9603 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2482 N$9724 N$9726 N$9605 N$9611 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2483 N$34849 N$9602 N$9613 N$9615 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2484 N$9608 N$34850 N$9617 N$9623 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2485 N$34851 N$9610 N$9625 N$9627 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2486 N$9612 N$34852 N$9629 N$9635 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2487 N$9614 N$9622 N$9637 N$34853 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2488 N$9620 N$9624 N$34854 N$9639 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2489 N$9626 N$9634 N$9641 N$34855 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2490 N$9632 N$9636 N$34856 N$9647 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2491 N$9638 N$9646 N$9774 N$9762 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2492 N$9644 N$9648 N$9764 N$9766 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2493 N$9604 N$9606 N$9607 N$9609 "Waveguide Crossing" sch_x=-4 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2494 N$9616 N$9618 N$9621 N$9619 "Waveguide Crossing" sch_x=0 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2495 N$9628 N$9630 N$9633 N$9631 "Waveguide Crossing" sch_x=0 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2496 N$9640 N$9642 N$9645 N$9643 "Waveguide Crossing" sch_x=4 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2497 N$9728 N$9730 N$9649 N$9651 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2498 N$9732 N$9736 N$9653 N$9659 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2499 N$34857 N$9650 N$9661 N$9663 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2500 N$9656 N$34858 N$9665 N$9671 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2501 N$34859 N$9658 N$9673 N$9675 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2502 N$9660 N$34860 N$9677 N$9683 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2503 N$9662 N$9670 N$9685 N$34861 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2504 N$9668 N$9672 N$34862 N$9687 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2505 N$9674 N$9682 N$9689 N$34863 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2506 N$9680 N$9684 N$34864 N$9695 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2507 N$9686 N$9694 N$9768 N$9770 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2508 N$9692 N$9696 N$9772 N$9776 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2509 N$9652 N$9654 N$9655 N$9657 "Waveguide Crossing" sch_x=-4 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2510 N$9664 N$9666 N$9669 N$9667 "Waveguide Crossing" sch_x=0 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2511 N$9676 N$9678 N$9681 N$9679 "Waveguide Crossing" sch_x=0 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2512 N$9688 N$9690 N$9693 N$9691 "Waveguide Crossing" sch_x=4 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2527 N$9761 N$9750 N$9737 N$9739 "Waveguide Crossing" sch_x=12 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2528 N$9752 N$9754 N$9741 N$9743 "Waveguide Crossing" sch_x=12 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2529 N$9756 N$9771 N$9745 N$9747 "Waveguide Crossing" sch_x=12 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2530 N$9763 N$9758 N$9749 N$9751 "Waveguide Crossing" sch_x=10 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2531 N$9760 N$9769 N$9753 N$9755 "Waveguide Crossing" sch_x=10 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2532 N$9765 N$9767 N$9757 N$9759 "Waveguide Crossing" sch_x=8 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2523 N$9773 N$9738 N$10238 N$10210 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2524 N$9740 N$9742 N$10212 N$10214 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2525 N$9744 N$9746 N$10216 N$10218 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2526 N$9748 N$9775 N$10220 N$10222 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2533 N$9910 N$9898 N$9777 N$9779 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2534 N$9900 N$9902 N$9781 N$9787 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2535 N$34865 N$9778 N$9789 N$9791 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2536 N$9784 N$34866 N$9793 N$9799 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2537 N$34867 N$9786 N$9801 N$9803 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2538 N$9788 N$34868 N$9805 N$9811 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2539 N$9790 N$9798 N$9813 N$34869 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2540 N$9796 N$9800 N$34870 N$9815 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2541 N$9802 N$9810 N$9817 N$34871 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2542 N$9808 N$9812 N$34872 N$9823 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2543 N$9814 N$9822 N$9950 N$9938 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2544 N$9820 N$9824 N$9940 N$9942 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2545 N$9780 N$9782 N$9783 N$9785 "Waveguide Crossing" sch_x=-4 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2546 N$9792 N$9794 N$9797 N$9795 "Waveguide Crossing" sch_x=0 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2547 N$9804 N$9806 N$9809 N$9807 "Waveguide Crossing" sch_x=0 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2548 N$9816 N$9818 N$9821 N$9819 "Waveguide Crossing" sch_x=4 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2549 N$9904 N$9906 N$9825 N$9827 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2550 N$9908 N$9912 N$9829 N$9835 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2551 N$34873 N$9826 N$9837 N$9839 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2552 N$9832 N$34874 N$9841 N$9847 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2553 N$34875 N$9834 N$9849 N$9851 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2554 N$9836 N$34876 N$9853 N$9859 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2555 N$9838 N$9846 N$9861 N$34877 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2556 N$9844 N$9848 N$34878 N$9863 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2557 N$9850 N$9858 N$9865 N$34879 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2558 N$9856 N$9860 N$34880 N$9871 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2559 N$9862 N$9870 N$9944 N$9946 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2560 N$9868 N$9872 N$9948 N$9952 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2561 N$9828 N$9830 N$9831 N$9833 "Waveguide Crossing" sch_x=-4 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2562 N$9840 N$9842 N$9845 N$9843 "Waveguide Crossing" sch_x=0 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2563 N$9852 N$9854 N$9857 N$9855 "Waveguide Crossing" sch_x=0 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2564 N$9864 N$9866 N$9869 N$9867 "Waveguide Crossing" sch_x=4 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2579 N$9937 N$9926 N$9913 N$9915 "Waveguide Crossing" sch_x=12 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2580 N$9928 N$9930 N$9917 N$9919 "Waveguide Crossing" sch_x=12 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2581 N$9932 N$9947 N$9921 N$9923 "Waveguide Crossing" sch_x=12 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2582 N$9939 N$9934 N$9925 N$9927 "Waveguide Crossing" sch_x=10 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2583 N$9936 N$9945 N$9929 N$9931 "Waveguide Crossing" sch_x=10 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2584 N$9941 N$9943 N$9933 N$9935 "Waveguide Crossing" sch_x=8 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2575 N$9949 N$9914 N$10224 N$10226 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2576 N$9916 N$9918 N$10228 N$10230 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2577 N$9920 N$9922 N$10232 N$10234 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2578 N$9924 N$9951 N$10236 N$10240 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2629 N$10209 N$10126 N$10097 N$10099 "Waveguide Crossing" sch_x=28 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2630 N$10128 N$10130 N$10101 N$10103 "Waveguide Crossing" sch_x=28 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2631 N$10132 N$10134 N$10105 N$10107 "Waveguide Crossing" sch_x=28 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2632 N$10136 N$10138 N$10109 N$10111 "Waveguide Crossing" sch_x=28 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2633 N$10140 N$10142 N$10113 N$10115 "Waveguide Crossing" sch_x=28 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2634 N$10144 N$10146 N$10117 N$10119 "Waveguide Crossing" sch_x=28 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2635 N$10148 N$10235 N$10121 N$10123 "Waveguide Crossing" sch_x=28 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2636 N$10211 N$10150 N$10125 N$10127 "Waveguide Crossing" sch_x=26 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2637 N$10152 N$10154 N$10129 N$10131 "Waveguide Crossing" sch_x=26 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2638 N$10156 N$10158 N$10133 N$10135 "Waveguide Crossing" sch_x=26 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2639 N$10160 N$10162 N$10137 N$10139 "Waveguide Crossing" sch_x=26 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2640 N$10164 N$10166 N$10141 N$10143 "Waveguide Crossing" sch_x=26 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2641 N$10168 N$10233 N$10145 N$10147 "Waveguide Crossing" sch_x=26 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2642 N$10213 N$10170 N$10149 N$10151 "Waveguide Crossing" sch_x=24 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2643 N$10172 N$10174 N$10153 N$10155 "Waveguide Crossing" sch_x=24 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2644 N$10176 N$10178 N$10157 N$10159 "Waveguide Crossing" sch_x=24 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2645 N$10180 N$10182 N$10161 N$10163 "Waveguide Crossing" sch_x=24 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2646 N$10184 N$10231 N$10165 N$10167 "Waveguide Crossing" sch_x=24 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2647 N$10215 N$10186 N$10169 N$10171 "Waveguide Crossing" sch_x=22 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2648 N$10188 N$10190 N$10173 N$10175 "Waveguide Crossing" sch_x=22 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2649 N$10192 N$10194 N$10177 N$10179 "Waveguide Crossing" sch_x=22 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2650 N$10196 N$10229 N$10181 N$10183 "Waveguide Crossing" sch_x=22 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2651 N$10217 N$10198 N$10185 N$10187 "Waveguide Crossing" sch_x=20 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2652 N$10200 N$10202 N$10189 N$10191 "Waveguide Crossing" sch_x=20 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2653 N$10204 N$10227 N$10193 N$10195 "Waveguide Crossing" sch_x=20 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2654 N$10219 N$10206 N$10197 N$10199 "Waveguide Crossing" sch_x=18 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2655 N$10208 N$10225 N$10201 N$10203 "Waveguide Crossing" sch_x=18 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2656 N$10221 N$10223 N$10205 N$10207 "Waveguide Crossing" sch_x=16 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2621 N$10237 N$10098 N$11296 N$11298 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2622 N$10100 N$10102 N$11300 N$11302 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2623 N$10104 N$10106 N$11304 N$11306 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2624 N$10108 N$10110 N$11308 N$11310 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2625 N$10112 N$10114 N$11312 N$11314 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2626 N$10116 N$10118 N$11316 N$11318 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2627 N$10120 N$10122 N$11320 N$11322 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2628 N$10124 N$10239 N$11324 N$11328 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2809 N$11265 N$10846 N$10785 N$10787 "Waveguide Crossing" sch_x=60 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2810 N$10848 N$10850 N$10789 N$10791 "Waveguide Crossing" sch_x=60 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2811 N$10852 N$10854 N$10793 N$10795 "Waveguide Crossing" sch_x=60 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2812 N$10856 N$10858 N$10797 N$10799 "Waveguide Crossing" sch_x=60 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2813 N$10860 N$10862 N$10801 N$10803 "Waveguide Crossing" sch_x=60 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2814 N$10864 N$10866 N$10805 N$10807 "Waveguide Crossing" sch_x=60 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2815 N$10868 N$10870 N$10809 N$10811 "Waveguide Crossing" sch_x=60 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2816 N$10872 N$10874 N$10813 N$10815 "Waveguide Crossing" sch_x=60 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2817 N$10876 N$10878 N$10817 N$10819 "Waveguide Crossing" sch_x=60 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2818 N$10880 N$10882 N$10821 N$10823 "Waveguide Crossing" sch_x=60 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2819 N$10884 N$10886 N$10825 N$10827 "Waveguide Crossing" sch_x=60 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2820 N$10888 N$10890 N$10829 N$10831 "Waveguide Crossing" sch_x=60 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2821 N$10892 N$10894 N$10833 N$10835 "Waveguide Crossing" sch_x=60 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2822 N$10896 N$10898 N$10837 N$10839 "Waveguide Crossing" sch_x=60 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2823 N$10900 N$11323 N$10841 N$10843 "Waveguide Crossing" sch_x=60 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2824 N$11267 N$10902 N$10845 N$10847 "Waveguide Crossing" sch_x=58 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2825 N$10904 N$10906 N$10849 N$10851 "Waveguide Crossing" sch_x=58 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2826 N$10908 N$10910 N$10853 N$10855 "Waveguide Crossing" sch_x=58 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2827 N$10912 N$10914 N$10857 N$10859 "Waveguide Crossing" sch_x=58 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2828 N$10916 N$10918 N$10861 N$10863 "Waveguide Crossing" sch_x=58 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2829 N$10920 N$10922 N$10865 N$10867 "Waveguide Crossing" sch_x=58 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2830 N$10924 N$10926 N$10869 N$10871 "Waveguide Crossing" sch_x=58 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2831 N$10928 N$10930 N$10873 N$10875 "Waveguide Crossing" sch_x=58 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2832 N$10932 N$10934 N$10877 N$10879 "Waveguide Crossing" sch_x=58 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2833 N$10936 N$10938 N$10881 N$10883 "Waveguide Crossing" sch_x=58 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2834 N$10940 N$10942 N$10885 N$10887 "Waveguide Crossing" sch_x=58 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2835 N$10944 N$10946 N$10889 N$10891 "Waveguide Crossing" sch_x=58 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2836 N$10948 N$10950 N$10893 N$10895 "Waveguide Crossing" sch_x=58 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2837 N$10952 N$11321 N$10897 N$10899 "Waveguide Crossing" sch_x=58 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2838 N$11269 N$10954 N$10901 N$10903 "Waveguide Crossing" sch_x=56 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2839 N$10956 N$10958 N$10905 N$10907 "Waveguide Crossing" sch_x=56 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2840 N$10960 N$10962 N$10909 N$10911 "Waveguide Crossing" sch_x=56 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2841 N$10964 N$10966 N$10913 N$10915 "Waveguide Crossing" sch_x=56 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2842 N$10968 N$10970 N$10917 N$10919 "Waveguide Crossing" sch_x=56 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2843 N$10972 N$10974 N$10921 N$10923 "Waveguide Crossing" sch_x=56 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2844 N$10976 N$10978 N$10925 N$10927 "Waveguide Crossing" sch_x=56 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2845 N$10980 N$10982 N$10929 N$10931 "Waveguide Crossing" sch_x=56 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2846 N$10984 N$10986 N$10933 N$10935 "Waveguide Crossing" sch_x=56 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2847 N$10988 N$10990 N$10937 N$10939 "Waveguide Crossing" sch_x=56 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2848 N$10992 N$10994 N$10941 N$10943 "Waveguide Crossing" sch_x=56 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2849 N$10996 N$10998 N$10945 N$10947 "Waveguide Crossing" sch_x=56 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2850 N$11000 N$11319 N$10949 N$10951 "Waveguide Crossing" sch_x=56 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2851 N$11271 N$11002 N$10953 N$10955 "Waveguide Crossing" sch_x=54 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2852 N$11004 N$11006 N$10957 N$10959 "Waveguide Crossing" sch_x=54 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2853 N$11008 N$11010 N$10961 N$10963 "Waveguide Crossing" sch_x=54 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2854 N$11012 N$11014 N$10965 N$10967 "Waveguide Crossing" sch_x=54 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2855 N$11016 N$11018 N$10969 N$10971 "Waveguide Crossing" sch_x=54 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2856 N$11020 N$11022 N$10973 N$10975 "Waveguide Crossing" sch_x=54 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2857 N$11024 N$11026 N$10977 N$10979 "Waveguide Crossing" sch_x=54 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2858 N$11028 N$11030 N$10981 N$10983 "Waveguide Crossing" sch_x=54 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2859 N$11032 N$11034 N$10985 N$10987 "Waveguide Crossing" sch_x=54 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2860 N$11036 N$11038 N$10989 N$10991 "Waveguide Crossing" sch_x=54 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2861 N$11040 N$11042 N$10993 N$10995 "Waveguide Crossing" sch_x=54 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2862 N$11044 N$11317 N$10997 N$10999 "Waveguide Crossing" sch_x=54 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2863 N$11273 N$11046 N$11001 N$11003 "Waveguide Crossing" sch_x=52 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2864 N$11048 N$11050 N$11005 N$11007 "Waveguide Crossing" sch_x=52 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2865 N$11052 N$11054 N$11009 N$11011 "Waveguide Crossing" sch_x=52 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2866 N$11056 N$11058 N$11013 N$11015 "Waveguide Crossing" sch_x=52 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2867 N$11060 N$11062 N$11017 N$11019 "Waveguide Crossing" sch_x=52 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2868 N$11064 N$11066 N$11021 N$11023 "Waveguide Crossing" sch_x=52 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2869 N$11068 N$11070 N$11025 N$11027 "Waveguide Crossing" sch_x=52 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2870 N$11072 N$11074 N$11029 N$11031 "Waveguide Crossing" sch_x=52 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2871 N$11076 N$11078 N$11033 N$11035 "Waveguide Crossing" sch_x=52 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2872 N$11080 N$11082 N$11037 N$11039 "Waveguide Crossing" sch_x=52 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2873 N$11084 N$11315 N$11041 N$11043 "Waveguide Crossing" sch_x=52 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2874 N$11275 N$11086 N$11045 N$11047 "Waveguide Crossing" sch_x=50 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2875 N$11088 N$11090 N$11049 N$11051 "Waveguide Crossing" sch_x=50 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2876 N$11092 N$11094 N$11053 N$11055 "Waveguide Crossing" sch_x=50 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2877 N$11096 N$11098 N$11057 N$11059 "Waveguide Crossing" sch_x=50 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2878 N$11100 N$11102 N$11061 N$11063 "Waveguide Crossing" sch_x=50 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2879 N$11104 N$11106 N$11065 N$11067 "Waveguide Crossing" sch_x=50 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2880 N$11108 N$11110 N$11069 N$11071 "Waveguide Crossing" sch_x=50 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2881 N$11112 N$11114 N$11073 N$11075 "Waveguide Crossing" sch_x=50 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2882 N$11116 N$11118 N$11077 N$11079 "Waveguide Crossing" sch_x=50 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2883 N$11120 N$11313 N$11081 N$11083 "Waveguide Crossing" sch_x=50 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2884 N$11277 N$11122 N$11085 N$11087 "Waveguide Crossing" sch_x=48 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2885 N$11124 N$11126 N$11089 N$11091 "Waveguide Crossing" sch_x=48 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2886 N$11128 N$11130 N$11093 N$11095 "Waveguide Crossing" sch_x=48 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2887 N$11132 N$11134 N$11097 N$11099 "Waveguide Crossing" sch_x=48 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2888 N$11136 N$11138 N$11101 N$11103 "Waveguide Crossing" sch_x=48 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2889 N$11140 N$11142 N$11105 N$11107 "Waveguide Crossing" sch_x=48 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2890 N$11144 N$11146 N$11109 N$11111 "Waveguide Crossing" sch_x=48 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2891 N$11148 N$11150 N$11113 N$11115 "Waveguide Crossing" sch_x=48 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2892 N$11152 N$11311 N$11117 N$11119 "Waveguide Crossing" sch_x=48 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2893 N$11279 N$11154 N$11121 N$11123 "Waveguide Crossing" sch_x=46 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2894 N$11156 N$11158 N$11125 N$11127 "Waveguide Crossing" sch_x=46 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2895 N$11160 N$11162 N$11129 N$11131 "Waveguide Crossing" sch_x=46 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2896 N$11164 N$11166 N$11133 N$11135 "Waveguide Crossing" sch_x=46 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2897 N$11168 N$11170 N$11137 N$11139 "Waveguide Crossing" sch_x=46 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2898 N$11172 N$11174 N$11141 N$11143 "Waveguide Crossing" sch_x=46 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2899 N$11176 N$11178 N$11145 N$11147 "Waveguide Crossing" sch_x=46 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2900 N$11180 N$11309 N$11149 N$11151 "Waveguide Crossing" sch_x=46 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2901 N$11281 N$11182 N$11153 N$11155 "Waveguide Crossing" sch_x=44 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2902 N$11184 N$11186 N$11157 N$11159 "Waveguide Crossing" sch_x=44 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2903 N$11188 N$11190 N$11161 N$11163 "Waveguide Crossing" sch_x=44 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2904 N$11192 N$11194 N$11165 N$11167 "Waveguide Crossing" sch_x=44 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2905 N$11196 N$11198 N$11169 N$11171 "Waveguide Crossing" sch_x=44 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2906 N$11200 N$11202 N$11173 N$11175 "Waveguide Crossing" sch_x=44 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2907 N$11204 N$11307 N$11177 N$11179 "Waveguide Crossing" sch_x=44 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2908 N$11283 N$11206 N$11181 N$11183 "Waveguide Crossing" sch_x=42 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2909 N$11208 N$11210 N$11185 N$11187 "Waveguide Crossing" sch_x=42 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2910 N$11212 N$11214 N$11189 N$11191 "Waveguide Crossing" sch_x=42 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2911 N$11216 N$11218 N$11193 N$11195 "Waveguide Crossing" sch_x=42 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2912 N$11220 N$11222 N$11197 N$11199 "Waveguide Crossing" sch_x=42 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2913 N$11224 N$11305 N$11201 N$11203 "Waveguide Crossing" sch_x=42 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2914 N$11285 N$11226 N$11205 N$11207 "Waveguide Crossing" sch_x=40 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2915 N$11228 N$11230 N$11209 N$11211 "Waveguide Crossing" sch_x=40 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2916 N$11232 N$11234 N$11213 N$11215 "Waveguide Crossing" sch_x=40 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2917 N$11236 N$11238 N$11217 N$11219 "Waveguide Crossing" sch_x=40 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2918 N$11240 N$11303 N$11221 N$11223 "Waveguide Crossing" sch_x=40 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2919 N$11287 N$11242 N$11225 N$11227 "Waveguide Crossing" sch_x=38 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2920 N$11244 N$11246 N$11229 N$11231 "Waveguide Crossing" sch_x=38 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2921 N$11248 N$11250 N$11233 N$11235 "Waveguide Crossing" sch_x=38 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2922 N$11252 N$11301 N$11237 N$11239 "Waveguide Crossing" sch_x=38 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2923 N$11289 N$11254 N$11241 N$11243 "Waveguide Crossing" sch_x=36 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2924 N$11256 N$11258 N$11245 N$11247 "Waveguide Crossing" sch_x=36 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2925 N$11260 N$11299 N$11249 N$11251 "Waveguide Crossing" sch_x=36 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2926 N$11291 N$11262 N$11253 N$11255 "Waveguide Crossing" sch_x=34 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2927 N$11264 N$11297 N$11257 N$11259 "Waveguide Crossing" sch_x=34 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2928 N$11293 N$11295 N$11261 N$11263 "Waveguide Crossing" sch_x=32 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2793 N$11325 N$10786 N$17918 N$17794 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2794 N$10788 N$10790 N$17796 N$17798 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2795 N$10792 N$10794 N$17800 N$17802 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2796 N$10796 N$10798 N$17804 N$17806 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2797 N$10800 N$10802 N$17808 N$17810 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2798 N$10804 N$10806 N$17812 N$17814 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2799 N$10808 N$10810 N$17816 N$17818 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2800 N$10812 N$10814 N$17820 N$17822 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2801 N$10816 N$10818 N$17824 N$17826 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2802 N$10820 N$10822 N$17828 N$17830 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2803 N$10824 N$10826 N$17832 N$17834 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2804 N$10828 N$10830 N$17836 N$17838 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2805 N$10832 N$10834 N$17840 N$17842 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2806 N$10836 N$10838 N$17844 N$17846 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2807 N$10840 N$10842 N$17848 N$17850 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2808 N$10844 N$11327 N$17852 N$17854 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2929 N$11462 N$11450 N$11329 N$11331 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-33.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2930 N$11452 N$11454 N$11333 N$11339 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-34.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2931 N$34881 N$11330 N$11341 N$11343 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2932 N$11336 N$34882 N$11345 N$11351 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2933 N$34883 N$11338 N$11353 N$11355 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2934 N$11340 N$34884 N$11357 N$11363 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2935 N$11342 N$11350 N$11365 N$34885 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2936 N$11348 N$11352 N$34886 N$11367 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2937 N$11354 N$11362 N$11369 N$34887 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2938 N$11360 N$11364 N$34888 N$11375 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2939 N$11366 N$11374 N$11502 N$11490 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-33.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2940 N$11372 N$11376 N$11492 N$11494 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-34.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2941 N$11332 N$11334 N$11335 N$11337 "Waveguide Crossing" sch_x=-4 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2942 N$11344 N$11346 N$11349 N$11347 "Waveguide Crossing" sch_x=0 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2943 N$11356 N$11358 N$11361 N$11359 "Waveguide Crossing" sch_x=0 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2944 N$11368 N$11370 N$11373 N$11371 "Waveguide Crossing" sch_x=4 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2945 N$11456 N$11458 N$11377 N$11379 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-37.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2946 N$11460 N$11464 N$11381 N$11387 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-38.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2947 N$34889 N$11378 N$11389 N$11391 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2948 N$11384 N$34890 N$11393 N$11399 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2949 N$34891 N$11386 N$11401 N$11403 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2950 N$11388 N$34892 N$11405 N$11411 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2951 N$11390 N$11398 N$11413 N$34893 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2952 N$11396 N$11400 N$34894 N$11415 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2953 N$11402 N$11410 N$11417 N$34895 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2954 N$11408 N$11412 N$34896 N$11423 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2955 N$11414 N$11422 N$11496 N$11498 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-37.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2956 N$11420 N$11424 N$11500 N$11504 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-38.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2957 N$11380 N$11382 N$11383 N$11385 "Waveguide Crossing" sch_x=-4 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2958 N$11392 N$11394 N$11397 N$11395 "Waveguide Crossing" sch_x=0 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2959 N$11404 N$11406 N$11409 N$11407 "Waveguide Crossing" sch_x=0 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2960 N$11416 N$11418 N$11421 N$11419 "Waveguide Crossing" sch_x=4 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2975 N$11489 N$11478 N$11465 N$11467 "Waveguide Crossing" sch_x=12 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2976 N$11480 N$11482 N$11469 N$11471 "Waveguide Crossing" sch_x=12 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2977 N$11484 N$11499 N$11473 N$11475 "Waveguide Crossing" sch_x=12 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2978 N$11491 N$11486 N$11477 N$11479 "Waveguide Crossing" sch_x=10 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2979 N$11488 N$11497 N$11481 N$11483 "Waveguide Crossing" sch_x=10 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2980 N$11493 N$11495 N$11485 N$11487 "Waveguide Crossing" sch_x=8 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2971 N$11501 N$11466 N$11966 N$11938 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2972 N$11468 N$11470 N$11940 N$11942 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2973 N$11472 N$11474 N$11944 N$11946 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2974 N$11476 N$11503 N$11948 N$11950 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2981 N$11638 N$11626 N$11505 N$11507 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-41.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2982 N$11628 N$11630 N$11509 N$11515 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-42.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2983 N$34897 N$11506 N$11517 N$11519 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2984 N$11512 N$34898 N$11521 N$11527 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2985 N$34899 N$11514 N$11529 N$11531 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2986 N$11516 N$34900 N$11533 N$11539 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2987 N$11518 N$11526 N$11541 N$34901 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2988 N$11524 N$11528 N$34902 N$11543 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2989 N$11530 N$11538 N$11545 N$34903 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2990 N$11536 N$11540 N$34904 N$11551 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2991 N$11542 N$11550 N$11678 N$11666 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-41.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2992 N$11548 N$11552 N$11668 N$11670 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-42.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2993 N$11508 N$11510 N$11511 N$11513 "Waveguide Crossing" sch_x=-4 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2994 N$11520 N$11522 N$11525 N$11523 "Waveguide Crossing" sch_x=0 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2995 N$11532 N$11534 N$11537 N$11535 "Waveguide Crossing" sch_x=0 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2996 N$11544 N$11546 N$11549 N$11547 "Waveguide Crossing" sch_x=4 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2997 N$11632 N$11634 N$11553 N$11555 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-45.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2998 N$11636 N$11640 N$11557 N$11563 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-46.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2999 N$34905 N$11554 N$11565 N$11567 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3000 N$11560 N$34906 N$11569 N$11575 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3001 N$34907 N$11562 N$11577 N$11579 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3002 N$11564 N$34908 N$11581 N$11587 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3003 N$11566 N$11574 N$11589 N$34909 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3004 N$11572 N$11576 N$34910 N$11591 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3005 N$11578 N$11586 N$11593 N$34911 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3006 N$11584 N$11588 N$34912 N$11599 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3007 N$11590 N$11598 N$11672 N$11674 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-45.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3008 N$11596 N$11600 N$11676 N$11680 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-46.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3009 N$11556 N$11558 N$11559 N$11561 "Waveguide Crossing" sch_x=-4 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3010 N$11568 N$11570 N$11573 N$11571 "Waveguide Crossing" sch_x=0 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3011 N$11580 N$11582 N$11585 N$11583 "Waveguide Crossing" sch_x=0 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3012 N$11592 N$11594 N$11597 N$11595 "Waveguide Crossing" sch_x=4 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3027 N$11665 N$11654 N$11641 N$11643 "Waveguide Crossing" sch_x=12 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3028 N$11656 N$11658 N$11645 N$11647 "Waveguide Crossing" sch_x=12 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3029 N$11660 N$11675 N$11649 N$11651 "Waveguide Crossing" sch_x=12 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3030 N$11667 N$11662 N$11653 N$11655 "Waveguide Crossing" sch_x=10 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3031 N$11664 N$11673 N$11657 N$11659 "Waveguide Crossing" sch_x=10 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3032 N$11669 N$11671 N$11661 N$11663 "Waveguide Crossing" sch_x=8 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3023 N$11677 N$11642 N$11952 N$11954 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3024 N$11644 N$11646 N$11956 N$11958 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3025 N$11648 N$11650 N$11960 N$11962 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3026 N$11652 N$11679 N$11964 N$11968 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3077 N$11937 N$11854 N$11825 N$11827 "Waveguide Crossing" sch_x=28 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3078 N$11856 N$11858 N$11829 N$11831 "Waveguide Crossing" sch_x=28 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3079 N$11860 N$11862 N$11833 N$11835 "Waveguide Crossing" sch_x=28 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3080 N$11864 N$11866 N$11837 N$11839 "Waveguide Crossing" sch_x=28 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3081 N$11868 N$11870 N$11841 N$11843 "Waveguide Crossing" sch_x=28 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3082 N$11872 N$11874 N$11845 N$11847 "Waveguide Crossing" sch_x=28 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3083 N$11876 N$11963 N$11849 N$11851 "Waveguide Crossing" sch_x=28 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3084 N$11939 N$11878 N$11853 N$11855 "Waveguide Crossing" sch_x=26 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3085 N$11880 N$11882 N$11857 N$11859 "Waveguide Crossing" sch_x=26 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3086 N$11884 N$11886 N$11861 N$11863 "Waveguide Crossing" sch_x=26 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3087 N$11888 N$11890 N$11865 N$11867 "Waveguide Crossing" sch_x=26 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3088 N$11892 N$11894 N$11869 N$11871 "Waveguide Crossing" sch_x=26 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3089 N$11896 N$11961 N$11873 N$11875 "Waveguide Crossing" sch_x=26 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3090 N$11941 N$11898 N$11877 N$11879 "Waveguide Crossing" sch_x=24 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3091 N$11900 N$11902 N$11881 N$11883 "Waveguide Crossing" sch_x=24 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3092 N$11904 N$11906 N$11885 N$11887 "Waveguide Crossing" sch_x=24 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3093 N$11908 N$11910 N$11889 N$11891 "Waveguide Crossing" sch_x=24 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3094 N$11912 N$11959 N$11893 N$11895 "Waveguide Crossing" sch_x=24 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3095 N$11943 N$11914 N$11897 N$11899 "Waveguide Crossing" sch_x=22 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3096 N$11916 N$11918 N$11901 N$11903 "Waveguide Crossing" sch_x=22 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3097 N$11920 N$11922 N$11905 N$11907 "Waveguide Crossing" sch_x=22 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3098 N$11924 N$11957 N$11909 N$11911 "Waveguide Crossing" sch_x=22 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3099 N$11945 N$11926 N$11913 N$11915 "Waveguide Crossing" sch_x=20 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3100 N$11928 N$11930 N$11917 N$11919 "Waveguide Crossing" sch_x=20 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3101 N$11932 N$11955 N$11921 N$11923 "Waveguide Crossing" sch_x=20 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3102 N$11947 N$11934 N$11925 N$11927 "Waveguide Crossing" sch_x=18 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3103 N$11936 N$11953 N$11929 N$11931 "Waveguide Crossing" sch_x=18 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3104 N$11949 N$11951 N$11933 N$11935 "Waveguide Crossing" sch_x=16 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3069 N$11965 N$11826 N$13694 N$13634 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3070 N$11828 N$11830 N$13636 N$13638 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3071 N$11832 N$11834 N$13640 N$13642 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3072 N$11836 N$11838 N$13644 N$13646 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3073 N$11840 N$11842 N$13648 N$13650 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3074 N$11844 N$11846 N$13652 N$13654 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3075 N$11848 N$11850 N$13656 N$13658 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3076 N$11852 N$11967 N$13660 N$13662 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3105 N$12102 N$12090 N$11969 N$11971 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-49.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3106 N$12092 N$12094 N$11973 N$11979 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-50.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3107 N$34913 N$11970 N$11981 N$11983 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3108 N$11976 N$34914 N$11985 N$11991 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3109 N$34915 N$11978 N$11993 N$11995 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3110 N$11980 N$34916 N$11997 N$12003 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3111 N$11982 N$11990 N$12005 N$34917 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3112 N$11988 N$11992 N$34918 N$12007 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3113 N$11994 N$12002 N$12009 N$34919 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3114 N$12000 N$12004 N$34920 N$12015 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3115 N$12006 N$12014 N$12142 N$12130 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-49.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3116 N$12012 N$12016 N$12132 N$12134 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-50.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3117 N$11972 N$11974 N$11975 N$11977 "Waveguide Crossing" sch_x=-4 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3118 N$11984 N$11986 N$11989 N$11987 "Waveguide Crossing" sch_x=0 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3119 N$11996 N$11998 N$12001 N$11999 "Waveguide Crossing" sch_x=0 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3120 N$12008 N$12010 N$12013 N$12011 "Waveguide Crossing" sch_x=4 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3121 N$12096 N$12098 N$12017 N$12019 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-53.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3122 N$12100 N$12104 N$12021 N$12027 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-54.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3123 N$34921 N$12018 N$12029 N$12031 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3124 N$12024 N$34922 N$12033 N$12039 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3125 N$34923 N$12026 N$12041 N$12043 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3126 N$12028 N$34924 N$12045 N$12051 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3127 N$12030 N$12038 N$12053 N$34925 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3128 N$12036 N$12040 N$34926 N$12055 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3129 N$12042 N$12050 N$12057 N$34927 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3130 N$12048 N$12052 N$34928 N$12063 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3131 N$12054 N$12062 N$12136 N$12138 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-53.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3132 N$12060 N$12064 N$12140 N$12144 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-54.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3133 N$12020 N$12022 N$12023 N$12025 "Waveguide Crossing" sch_x=-4 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3134 N$12032 N$12034 N$12037 N$12035 "Waveguide Crossing" sch_x=0 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3135 N$12044 N$12046 N$12049 N$12047 "Waveguide Crossing" sch_x=0 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3136 N$12056 N$12058 N$12061 N$12059 "Waveguide Crossing" sch_x=4 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3151 N$12129 N$12118 N$12105 N$12107 "Waveguide Crossing" sch_x=12 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3152 N$12120 N$12122 N$12109 N$12111 "Waveguide Crossing" sch_x=12 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3153 N$12124 N$12139 N$12113 N$12115 "Waveguide Crossing" sch_x=12 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3154 N$12131 N$12126 N$12117 N$12119 "Waveguide Crossing" sch_x=10 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3155 N$12128 N$12137 N$12121 N$12123 "Waveguide Crossing" sch_x=10 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3156 N$12133 N$12135 N$12125 N$12127 "Waveguide Crossing" sch_x=8 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3147 N$12141 N$12106 N$12606 N$12578 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3148 N$12108 N$12110 N$12580 N$12582 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3149 N$12112 N$12114 N$12584 N$12586 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3150 N$12116 N$12143 N$12588 N$12590 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3157 N$12278 N$12266 N$12145 N$12147 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-57.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3158 N$12268 N$12270 N$12149 N$12155 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-58.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3159 N$34929 N$12146 N$12157 N$12159 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3160 N$12152 N$34930 N$12161 N$12167 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3161 N$34931 N$12154 N$12169 N$12171 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3162 N$12156 N$34932 N$12173 N$12179 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3163 N$12158 N$12166 N$12181 N$34933 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3164 N$12164 N$12168 N$34934 N$12183 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3165 N$12170 N$12178 N$12185 N$34935 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3166 N$12176 N$12180 N$34936 N$12191 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3167 N$12182 N$12190 N$12318 N$12306 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-57.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3168 N$12188 N$12192 N$12308 N$12310 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-58.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3169 N$12148 N$12150 N$12151 N$12153 "Waveguide Crossing" sch_x=-4 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3170 N$12160 N$12162 N$12165 N$12163 "Waveguide Crossing" sch_x=0 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3171 N$12172 N$12174 N$12177 N$12175 "Waveguide Crossing" sch_x=0 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3172 N$12184 N$12186 N$12189 N$12187 "Waveguide Crossing" sch_x=4 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3173 N$12272 N$12274 N$12193 N$12195 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-61.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3174 N$12276 N$12280 N$12197 N$12203 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-62.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3175 N$34937 N$12194 N$12205 N$12207 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3176 N$12200 N$34938 N$12209 N$12215 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3177 N$34939 N$12202 N$12217 N$12219 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3178 N$12204 N$34940 N$12221 N$12227 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-63.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3179 N$12206 N$12214 N$12229 N$34941 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3180 N$12212 N$12216 N$34942 N$12231 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3181 N$12218 N$12226 N$12233 N$34943 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3182 N$12224 N$12228 N$34944 N$12239 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-63.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3183 N$12230 N$12238 N$12312 N$12314 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-61.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3184 N$12236 N$12240 N$12316 N$12320 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-62.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3185 N$12196 N$12198 N$12199 N$12201 "Waveguide Crossing" sch_x=-4 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3186 N$12208 N$12210 N$12213 N$12211 "Waveguide Crossing" sch_x=0 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3187 N$12220 N$12222 N$12225 N$12223 "Waveguide Crossing" sch_x=0 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3188 N$12232 N$12234 N$12237 N$12235 "Waveguide Crossing" sch_x=4 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3203 N$12305 N$12294 N$12281 N$12283 "Waveguide Crossing" sch_x=12 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3204 N$12296 N$12298 N$12285 N$12287 "Waveguide Crossing" sch_x=12 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3205 N$12300 N$12315 N$12289 N$12291 "Waveguide Crossing" sch_x=12 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3206 N$12307 N$12302 N$12293 N$12295 "Waveguide Crossing" sch_x=10 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3207 N$12304 N$12313 N$12297 N$12299 "Waveguide Crossing" sch_x=10 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3208 N$12309 N$12311 N$12301 N$12303 "Waveguide Crossing" sch_x=8 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3199 N$12317 N$12282 N$12592 N$12594 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3200 N$12284 N$12286 N$12596 N$12598 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3201 N$12288 N$12290 N$12600 N$12602 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3202 N$12292 N$12319 N$12604 N$12608 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3253 N$12577 N$12494 N$12465 N$12467 "Waveguide Crossing" sch_x=28 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3254 N$12496 N$12498 N$12469 N$12471 "Waveguide Crossing" sch_x=28 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3255 N$12500 N$12502 N$12473 N$12475 "Waveguide Crossing" sch_x=28 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3256 N$12504 N$12506 N$12477 N$12479 "Waveguide Crossing" sch_x=28 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3257 N$12508 N$12510 N$12481 N$12483 "Waveguide Crossing" sch_x=28 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3258 N$12512 N$12514 N$12485 N$12487 "Waveguide Crossing" sch_x=28 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3259 N$12516 N$12603 N$12489 N$12491 "Waveguide Crossing" sch_x=28 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3260 N$12579 N$12518 N$12493 N$12495 "Waveguide Crossing" sch_x=26 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3261 N$12520 N$12522 N$12497 N$12499 "Waveguide Crossing" sch_x=26 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3262 N$12524 N$12526 N$12501 N$12503 "Waveguide Crossing" sch_x=26 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3263 N$12528 N$12530 N$12505 N$12507 "Waveguide Crossing" sch_x=26 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3264 N$12532 N$12534 N$12509 N$12511 "Waveguide Crossing" sch_x=26 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3265 N$12536 N$12601 N$12513 N$12515 "Waveguide Crossing" sch_x=26 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3266 N$12581 N$12538 N$12517 N$12519 "Waveguide Crossing" sch_x=24 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3267 N$12540 N$12542 N$12521 N$12523 "Waveguide Crossing" sch_x=24 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3268 N$12544 N$12546 N$12525 N$12527 "Waveguide Crossing" sch_x=24 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3269 N$12548 N$12550 N$12529 N$12531 "Waveguide Crossing" sch_x=24 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3270 N$12552 N$12599 N$12533 N$12535 "Waveguide Crossing" sch_x=24 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3271 N$12583 N$12554 N$12537 N$12539 "Waveguide Crossing" sch_x=22 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3272 N$12556 N$12558 N$12541 N$12543 "Waveguide Crossing" sch_x=22 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3273 N$12560 N$12562 N$12545 N$12547 "Waveguide Crossing" sch_x=22 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3274 N$12564 N$12597 N$12549 N$12551 "Waveguide Crossing" sch_x=22 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3275 N$12585 N$12566 N$12553 N$12555 "Waveguide Crossing" sch_x=20 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3276 N$12568 N$12570 N$12557 N$12559 "Waveguide Crossing" sch_x=20 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3277 N$12572 N$12595 N$12561 N$12563 "Waveguide Crossing" sch_x=20 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3278 N$12587 N$12574 N$12565 N$12567 "Waveguide Crossing" sch_x=18 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3279 N$12576 N$12593 N$12569 N$12571 "Waveguide Crossing" sch_x=18 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3280 N$12589 N$12591 N$12573 N$12575 "Waveguide Crossing" sch_x=16 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3245 N$12605 N$12466 N$13664 N$13666 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3246 N$12468 N$12470 N$13668 N$13670 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3247 N$12472 N$12474 N$13672 N$13674 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3248 N$12476 N$12478 N$13676 N$13678 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3249 N$12480 N$12482 N$13680 N$13682 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3250 N$12484 N$12486 N$13684 N$13686 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3251 N$12488 N$12490 N$13688 N$13690 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3252 N$12492 N$12607 N$13692 N$13696 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3433 N$13633 N$13214 N$13153 N$13155 "Waveguide Crossing" sch_x=60 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3434 N$13216 N$13218 N$13157 N$13159 "Waveguide Crossing" sch_x=60 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3435 N$13220 N$13222 N$13161 N$13163 "Waveguide Crossing" sch_x=60 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3436 N$13224 N$13226 N$13165 N$13167 "Waveguide Crossing" sch_x=60 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3437 N$13228 N$13230 N$13169 N$13171 "Waveguide Crossing" sch_x=60 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3438 N$13232 N$13234 N$13173 N$13175 "Waveguide Crossing" sch_x=60 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3439 N$13236 N$13238 N$13177 N$13179 "Waveguide Crossing" sch_x=60 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3440 N$13240 N$13242 N$13181 N$13183 "Waveguide Crossing" sch_x=60 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3441 N$13244 N$13246 N$13185 N$13187 "Waveguide Crossing" sch_x=60 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3442 N$13248 N$13250 N$13189 N$13191 "Waveguide Crossing" sch_x=60 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3443 N$13252 N$13254 N$13193 N$13195 "Waveguide Crossing" sch_x=60 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3444 N$13256 N$13258 N$13197 N$13199 "Waveguide Crossing" sch_x=60 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3445 N$13260 N$13262 N$13201 N$13203 "Waveguide Crossing" sch_x=60 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3446 N$13264 N$13266 N$13205 N$13207 "Waveguide Crossing" sch_x=60 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3447 N$13268 N$13691 N$13209 N$13211 "Waveguide Crossing" sch_x=60 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3448 N$13635 N$13270 N$13213 N$13215 "Waveguide Crossing" sch_x=58 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3449 N$13272 N$13274 N$13217 N$13219 "Waveguide Crossing" sch_x=58 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3450 N$13276 N$13278 N$13221 N$13223 "Waveguide Crossing" sch_x=58 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3451 N$13280 N$13282 N$13225 N$13227 "Waveguide Crossing" sch_x=58 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3452 N$13284 N$13286 N$13229 N$13231 "Waveguide Crossing" sch_x=58 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3453 N$13288 N$13290 N$13233 N$13235 "Waveguide Crossing" sch_x=58 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3454 N$13292 N$13294 N$13237 N$13239 "Waveguide Crossing" sch_x=58 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3455 N$13296 N$13298 N$13241 N$13243 "Waveguide Crossing" sch_x=58 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3456 N$13300 N$13302 N$13245 N$13247 "Waveguide Crossing" sch_x=58 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3457 N$13304 N$13306 N$13249 N$13251 "Waveguide Crossing" sch_x=58 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3458 N$13308 N$13310 N$13253 N$13255 "Waveguide Crossing" sch_x=58 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3459 N$13312 N$13314 N$13257 N$13259 "Waveguide Crossing" sch_x=58 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3460 N$13316 N$13318 N$13261 N$13263 "Waveguide Crossing" sch_x=58 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3461 N$13320 N$13689 N$13265 N$13267 "Waveguide Crossing" sch_x=58 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3462 N$13637 N$13322 N$13269 N$13271 "Waveguide Crossing" sch_x=56 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3463 N$13324 N$13326 N$13273 N$13275 "Waveguide Crossing" sch_x=56 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3464 N$13328 N$13330 N$13277 N$13279 "Waveguide Crossing" sch_x=56 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3465 N$13332 N$13334 N$13281 N$13283 "Waveguide Crossing" sch_x=56 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3466 N$13336 N$13338 N$13285 N$13287 "Waveguide Crossing" sch_x=56 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3467 N$13340 N$13342 N$13289 N$13291 "Waveguide Crossing" sch_x=56 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3468 N$13344 N$13346 N$13293 N$13295 "Waveguide Crossing" sch_x=56 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3469 N$13348 N$13350 N$13297 N$13299 "Waveguide Crossing" sch_x=56 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3470 N$13352 N$13354 N$13301 N$13303 "Waveguide Crossing" sch_x=56 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3471 N$13356 N$13358 N$13305 N$13307 "Waveguide Crossing" sch_x=56 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3472 N$13360 N$13362 N$13309 N$13311 "Waveguide Crossing" sch_x=56 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3473 N$13364 N$13366 N$13313 N$13315 "Waveguide Crossing" sch_x=56 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3474 N$13368 N$13687 N$13317 N$13319 "Waveguide Crossing" sch_x=56 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3475 N$13639 N$13370 N$13321 N$13323 "Waveguide Crossing" sch_x=54 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3476 N$13372 N$13374 N$13325 N$13327 "Waveguide Crossing" sch_x=54 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3477 N$13376 N$13378 N$13329 N$13331 "Waveguide Crossing" sch_x=54 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3478 N$13380 N$13382 N$13333 N$13335 "Waveguide Crossing" sch_x=54 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3479 N$13384 N$13386 N$13337 N$13339 "Waveguide Crossing" sch_x=54 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3480 N$13388 N$13390 N$13341 N$13343 "Waveguide Crossing" sch_x=54 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3481 N$13392 N$13394 N$13345 N$13347 "Waveguide Crossing" sch_x=54 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3482 N$13396 N$13398 N$13349 N$13351 "Waveguide Crossing" sch_x=54 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3483 N$13400 N$13402 N$13353 N$13355 "Waveguide Crossing" sch_x=54 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3484 N$13404 N$13406 N$13357 N$13359 "Waveguide Crossing" sch_x=54 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3485 N$13408 N$13410 N$13361 N$13363 "Waveguide Crossing" sch_x=54 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3486 N$13412 N$13685 N$13365 N$13367 "Waveguide Crossing" sch_x=54 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3487 N$13641 N$13414 N$13369 N$13371 "Waveguide Crossing" sch_x=52 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3488 N$13416 N$13418 N$13373 N$13375 "Waveguide Crossing" sch_x=52 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3489 N$13420 N$13422 N$13377 N$13379 "Waveguide Crossing" sch_x=52 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3490 N$13424 N$13426 N$13381 N$13383 "Waveguide Crossing" sch_x=52 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3491 N$13428 N$13430 N$13385 N$13387 "Waveguide Crossing" sch_x=52 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3492 N$13432 N$13434 N$13389 N$13391 "Waveguide Crossing" sch_x=52 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3493 N$13436 N$13438 N$13393 N$13395 "Waveguide Crossing" sch_x=52 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3494 N$13440 N$13442 N$13397 N$13399 "Waveguide Crossing" sch_x=52 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3495 N$13444 N$13446 N$13401 N$13403 "Waveguide Crossing" sch_x=52 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3496 N$13448 N$13450 N$13405 N$13407 "Waveguide Crossing" sch_x=52 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3497 N$13452 N$13683 N$13409 N$13411 "Waveguide Crossing" sch_x=52 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3498 N$13643 N$13454 N$13413 N$13415 "Waveguide Crossing" sch_x=50 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3499 N$13456 N$13458 N$13417 N$13419 "Waveguide Crossing" sch_x=50 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3500 N$13460 N$13462 N$13421 N$13423 "Waveguide Crossing" sch_x=50 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3501 N$13464 N$13466 N$13425 N$13427 "Waveguide Crossing" sch_x=50 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3502 N$13468 N$13470 N$13429 N$13431 "Waveguide Crossing" sch_x=50 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3503 N$13472 N$13474 N$13433 N$13435 "Waveguide Crossing" sch_x=50 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3504 N$13476 N$13478 N$13437 N$13439 "Waveguide Crossing" sch_x=50 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3505 N$13480 N$13482 N$13441 N$13443 "Waveguide Crossing" sch_x=50 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3506 N$13484 N$13486 N$13445 N$13447 "Waveguide Crossing" sch_x=50 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3507 N$13488 N$13681 N$13449 N$13451 "Waveguide Crossing" sch_x=50 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3508 N$13645 N$13490 N$13453 N$13455 "Waveguide Crossing" sch_x=48 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3509 N$13492 N$13494 N$13457 N$13459 "Waveguide Crossing" sch_x=48 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3510 N$13496 N$13498 N$13461 N$13463 "Waveguide Crossing" sch_x=48 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3511 N$13500 N$13502 N$13465 N$13467 "Waveguide Crossing" sch_x=48 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3512 N$13504 N$13506 N$13469 N$13471 "Waveguide Crossing" sch_x=48 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3513 N$13508 N$13510 N$13473 N$13475 "Waveguide Crossing" sch_x=48 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3514 N$13512 N$13514 N$13477 N$13479 "Waveguide Crossing" sch_x=48 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3515 N$13516 N$13518 N$13481 N$13483 "Waveguide Crossing" sch_x=48 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3516 N$13520 N$13679 N$13485 N$13487 "Waveguide Crossing" sch_x=48 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3517 N$13647 N$13522 N$13489 N$13491 "Waveguide Crossing" sch_x=46 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3518 N$13524 N$13526 N$13493 N$13495 "Waveguide Crossing" sch_x=46 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3519 N$13528 N$13530 N$13497 N$13499 "Waveguide Crossing" sch_x=46 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3520 N$13532 N$13534 N$13501 N$13503 "Waveguide Crossing" sch_x=46 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3521 N$13536 N$13538 N$13505 N$13507 "Waveguide Crossing" sch_x=46 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3522 N$13540 N$13542 N$13509 N$13511 "Waveguide Crossing" sch_x=46 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3523 N$13544 N$13546 N$13513 N$13515 "Waveguide Crossing" sch_x=46 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3524 N$13548 N$13677 N$13517 N$13519 "Waveguide Crossing" sch_x=46 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3525 N$13649 N$13550 N$13521 N$13523 "Waveguide Crossing" sch_x=44 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3526 N$13552 N$13554 N$13525 N$13527 "Waveguide Crossing" sch_x=44 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3527 N$13556 N$13558 N$13529 N$13531 "Waveguide Crossing" sch_x=44 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3528 N$13560 N$13562 N$13533 N$13535 "Waveguide Crossing" sch_x=44 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3529 N$13564 N$13566 N$13537 N$13539 "Waveguide Crossing" sch_x=44 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3530 N$13568 N$13570 N$13541 N$13543 "Waveguide Crossing" sch_x=44 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3531 N$13572 N$13675 N$13545 N$13547 "Waveguide Crossing" sch_x=44 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3532 N$13651 N$13574 N$13549 N$13551 "Waveguide Crossing" sch_x=42 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3533 N$13576 N$13578 N$13553 N$13555 "Waveguide Crossing" sch_x=42 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3534 N$13580 N$13582 N$13557 N$13559 "Waveguide Crossing" sch_x=42 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3535 N$13584 N$13586 N$13561 N$13563 "Waveguide Crossing" sch_x=42 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3536 N$13588 N$13590 N$13565 N$13567 "Waveguide Crossing" sch_x=42 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3537 N$13592 N$13673 N$13569 N$13571 "Waveguide Crossing" sch_x=42 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3538 N$13653 N$13594 N$13573 N$13575 "Waveguide Crossing" sch_x=40 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3539 N$13596 N$13598 N$13577 N$13579 "Waveguide Crossing" sch_x=40 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3540 N$13600 N$13602 N$13581 N$13583 "Waveguide Crossing" sch_x=40 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3541 N$13604 N$13606 N$13585 N$13587 "Waveguide Crossing" sch_x=40 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3542 N$13608 N$13671 N$13589 N$13591 "Waveguide Crossing" sch_x=40 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3543 N$13655 N$13610 N$13593 N$13595 "Waveguide Crossing" sch_x=38 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3544 N$13612 N$13614 N$13597 N$13599 "Waveguide Crossing" sch_x=38 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3545 N$13616 N$13618 N$13601 N$13603 "Waveguide Crossing" sch_x=38 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3546 N$13620 N$13669 N$13605 N$13607 "Waveguide Crossing" sch_x=38 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3547 N$13657 N$13622 N$13609 N$13611 "Waveguide Crossing" sch_x=36 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3548 N$13624 N$13626 N$13613 N$13615 "Waveguide Crossing" sch_x=36 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3549 N$13628 N$13667 N$13617 N$13619 "Waveguide Crossing" sch_x=36 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3550 N$13659 N$13630 N$13621 N$13623 "Waveguide Crossing" sch_x=34 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3551 N$13632 N$13665 N$13625 N$13627 "Waveguide Crossing" sch_x=34 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C3552 N$13661 N$13663 N$13629 N$13631 "Waveguide Crossing" sch_x=32 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3417 N$13693 N$13154 N$17856 N$17858 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3418 N$13156 N$13158 N$17860 N$17862 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3419 N$13160 N$13162 N$17864 N$17866 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3420 N$13164 N$13166 N$17868 N$17870 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3421 N$13168 N$13170 N$17872 N$17874 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3422 N$13172 N$13174 N$17876 N$17878 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3423 N$13176 N$13178 N$17880 N$17882 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3424 N$13180 N$13182 N$17884 N$17886 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3425 N$13184 N$13186 N$17888 N$17890 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3426 N$13188 N$13190 N$17892 N$17894 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3427 N$13192 N$13194 N$17896 N$17898 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3428 N$13196 N$13198 N$17900 N$17902 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3429 N$13200 N$13202 N$17904 N$17906 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3430 N$13204 N$13206 N$17908 N$17910 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3431 N$13208 N$13210 N$17912 N$17914 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3432 N$13212 N$13695 N$17916 N$17920 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4113 N$17793 N$15934 N$15809 N$15811 "Waveguide Crossing" sch_x=124 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4114 N$15936 N$15938 N$15813 N$15815 "Waveguide Crossing" sch_x=124 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4115 N$15940 N$15942 N$15817 N$15819 "Waveguide Crossing" sch_x=124 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4116 N$15944 N$15946 N$15821 N$15823 "Waveguide Crossing" sch_x=124 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4117 N$15948 N$15950 N$15825 N$15827 "Waveguide Crossing" sch_x=124 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4118 N$15952 N$15954 N$15829 N$15831 "Waveguide Crossing" sch_x=124 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4119 N$15956 N$15958 N$15833 N$15835 "Waveguide Crossing" sch_x=124 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4120 N$15960 N$15962 N$15837 N$15839 "Waveguide Crossing" sch_x=124 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4121 N$15964 N$15966 N$15841 N$15843 "Waveguide Crossing" sch_x=124 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4122 N$15968 N$15970 N$15845 N$15847 "Waveguide Crossing" sch_x=124 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4123 N$15972 N$15974 N$15849 N$15851 "Waveguide Crossing" sch_x=124 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4124 N$15976 N$15978 N$15853 N$15855 "Waveguide Crossing" sch_x=124 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4125 N$15980 N$15982 N$15857 N$15859 "Waveguide Crossing" sch_x=124 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4126 N$15984 N$15986 N$15861 N$15863 "Waveguide Crossing" sch_x=124 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4127 N$15988 N$15990 N$15865 N$15867 "Waveguide Crossing" sch_x=124 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4128 N$15992 N$15994 N$15869 N$15871 "Waveguide Crossing" sch_x=124 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4129 N$15996 N$15998 N$15873 N$15875 "Waveguide Crossing" sch_x=124 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4130 N$16000 N$16002 N$15877 N$15879 "Waveguide Crossing" sch_x=124 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4131 N$16004 N$16006 N$15881 N$15883 "Waveguide Crossing" sch_x=124 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4132 N$16008 N$16010 N$15885 N$15887 "Waveguide Crossing" sch_x=124 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4133 N$16012 N$16014 N$15889 N$15891 "Waveguide Crossing" sch_x=124 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4134 N$16016 N$16018 N$15893 N$15895 "Waveguide Crossing" sch_x=124 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4135 N$16020 N$16022 N$15897 N$15899 "Waveguide Crossing" sch_x=124 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4136 N$16024 N$16026 N$15901 N$15903 "Waveguide Crossing" sch_x=124 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4137 N$16028 N$16030 N$15905 N$15907 "Waveguide Crossing" sch_x=124 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4138 N$16032 N$16034 N$15909 N$15911 "Waveguide Crossing" sch_x=124 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4139 N$16036 N$16038 N$15913 N$15915 "Waveguide Crossing" sch_x=124 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4140 N$16040 N$16042 N$15917 N$15919 "Waveguide Crossing" sch_x=124 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4141 N$16044 N$16046 N$15921 N$15923 "Waveguide Crossing" sch_x=124 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4142 N$16048 N$16050 N$15925 N$15927 "Waveguide Crossing" sch_x=124 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4143 N$16052 N$17915 N$15929 N$15931 "Waveguide Crossing" sch_x=124 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4144 N$17795 N$16054 N$15933 N$15935 "Waveguide Crossing" sch_x=122 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4145 N$16056 N$16058 N$15937 N$15939 "Waveguide Crossing" sch_x=122 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4146 N$16060 N$16062 N$15941 N$15943 "Waveguide Crossing" sch_x=122 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4147 N$16064 N$16066 N$15945 N$15947 "Waveguide Crossing" sch_x=122 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4148 N$16068 N$16070 N$15949 N$15951 "Waveguide Crossing" sch_x=122 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4149 N$16072 N$16074 N$15953 N$15955 "Waveguide Crossing" sch_x=122 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4150 N$16076 N$16078 N$15957 N$15959 "Waveguide Crossing" sch_x=122 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4151 N$16080 N$16082 N$15961 N$15963 "Waveguide Crossing" sch_x=122 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4152 N$16084 N$16086 N$15965 N$15967 "Waveguide Crossing" sch_x=122 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4153 N$16088 N$16090 N$15969 N$15971 "Waveguide Crossing" sch_x=122 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4154 N$16092 N$16094 N$15973 N$15975 "Waveguide Crossing" sch_x=122 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4155 N$16096 N$16098 N$15977 N$15979 "Waveguide Crossing" sch_x=122 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4156 N$16100 N$16102 N$15981 N$15983 "Waveguide Crossing" sch_x=122 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4157 N$16104 N$16106 N$15985 N$15987 "Waveguide Crossing" sch_x=122 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4158 N$16108 N$16110 N$15989 N$15991 "Waveguide Crossing" sch_x=122 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4159 N$16112 N$16114 N$15993 N$15995 "Waveguide Crossing" sch_x=122 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4160 N$16116 N$16118 N$15997 N$15999 "Waveguide Crossing" sch_x=122 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4161 N$16120 N$16122 N$16001 N$16003 "Waveguide Crossing" sch_x=122 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4162 N$16124 N$16126 N$16005 N$16007 "Waveguide Crossing" sch_x=122 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4163 N$16128 N$16130 N$16009 N$16011 "Waveguide Crossing" sch_x=122 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4164 N$16132 N$16134 N$16013 N$16015 "Waveguide Crossing" sch_x=122 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4165 N$16136 N$16138 N$16017 N$16019 "Waveguide Crossing" sch_x=122 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4166 N$16140 N$16142 N$16021 N$16023 "Waveguide Crossing" sch_x=122 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4167 N$16144 N$16146 N$16025 N$16027 "Waveguide Crossing" sch_x=122 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4168 N$16148 N$16150 N$16029 N$16031 "Waveguide Crossing" sch_x=122 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4169 N$16152 N$16154 N$16033 N$16035 "Waveguide Crossing" sch_x=122 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4170 N$16156 N$16158 N$16037 N$16039 "Waveguide Crossing" sch_x=122 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4171 N$16160 N$16162 N$16041 N$16043 "Waveguide Crossing" sch_x=122 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4172 N$16164 N$16166 N$16045 N$16047 "Waveguide Crossing" sch_x=122 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4173 N$16168 N$17913 N$16049 N$16051 "Waveguide Crossing" sch_x=122 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4174 N$17797 N$16170 N$16053 N$16055 "Waveguide Crossing" sch_x=120 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4175 N$16172 N$16174 N$16057 N$16059 "Waveguide Crossing" sch_x=120 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4176 N$16176 N$16178 N$16061 N$16063 "Waveguide Crossing" sch_x=120 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4177 N$16180 N$16182 N$16065 N$16067 "Waveguide Crossing" sch_x=120 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4178 N$16184 N$16186 N$16069 N$16071 "Waveguide Crossing" sch_x=120 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4179 N$16188 N$16190 N$16073 N$16075 "Waveguide Crossing" sch_x=120 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4180 N$16192 N$16194 N$16077 N$16079 "Waveguide Crossing" sch_x=120 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4181 N$16196 N$16198 N$16081 N$16083 "Waveguide Crossing" sch_x=120 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4182 N$16200 N$16202 N$16085 N$16087 "Waveguide Crossing" sch_x=120 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4183 N$16204 N$16206 N$16089 N$16091 "Waveguide Crossing" sch_x=120 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4184 N$16208 N$16210 N$16093 N$16095 "Waveguide Crossing" sch_x=120 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4185 N$16212 N$16214 N$16097 N$16099 "Waveguide Crossing" sch_x=120 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4186 N$16216 N$16218 N$16101 N$16103 "Waveguide Crossing" sch_x=120 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4187 N$16220 N$16222 N$16105 N$16107 "Waveguide Crossing" sch_x=120 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4188 N$16224 N$16226 N$16109 N$16111 "Waveguide Crossing" sch_x=120 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4189 N$16228 N$16230 N$16113 N$16115 "Waveguide Crossing" sch_x=120 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4190 N$16232 N$16234 N$16117 N$16119 "Waveguide Crossing" sch_x=120 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4191 N$16236 N$16238 N$16121 N$16123 "Waveguide Crossing" sch_x=120 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4192 N$16240 N$16242 N$16125 N$16127 "Waveguide Crossing" sch_x=120 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4193 N$16244 N$16246 N$16129 N$16131 "Waveguide Crossing" sch_x=120 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4194 N$16248 N$16250 N$16133 N$16135 "Waveguide Crossing" sch_x=120 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4195 N$16252 N$16254 N$16137 N$16139 "Waveguide Crossing" sch_x=120 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4196 N$16256 N$16258 N$16141 N$16143 "Waveguide Crossing" sch_x=120 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4197 N$16260 N$16262 N$16145 N$16147 "Waveguide Crossing" sch_x=120 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4198 N$16264 N$16266 N$16149 N$16151 "Waveguide Crossing" sch_x=120 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4199 N$16268 N$16270 N$16153 N$16155 "Waveguide Crossing" sch_x=120 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4200 N$16272 N$16274 N$16157 N$16159 "Waveguide Crossing" sch_x=120 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4201 N$16276 N$16278 N$16161 N$16163 "Waveguide Crossing" sch_x=120 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4202 N$16280 N$17911 N$16165 N$16167 "Waveguide Crossing" sch_x=120 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4203 N$17799 N$16282 N$16169 N$16171 "Waveguide Crossing" sch_x=118 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4204 N$16284 N$16286 N$16173 N$16175 "Waveguide Crossing" sch_x=118 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4205 N$16288 N$16290 N$16177 N$16179 "Waveguide Crossing" sch_x=118 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4206 N$16292 N$16294 N$16181 N$16183 "Waveguide Crossing" sch_x=118 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4207 N$16296 N$16298 N$16185 N$16187 "Waveguide Crossing" sch_x=118 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4208 N$16300 N$16302 N$16189 N$16191 "Waveguide Crossing" sch_x=118 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4209 N$16304 N$16306 N$16193 N$16195 "Waveguide Crossing" sch_x=118 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4210 N$16308 N$16310 N$16197 N$16199 "Waveguide Crossing" sch_x=118 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4211 N$16312 N$16314 N$16201 N$16203 "Waveguide Crossing" sch_x=118 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4212 N$16316 N$16318 N$16205 N$16207 "Waveguide Crossing" sch_x=118 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4213 N$16320 N$16322 N$16209 N$16211 "Waveguide Crossing" sch_x=118 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4214 N$16324 N$16326 N$16213 N$16215 "Waveguide Crossing" sch_x=118 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4215 N$16328 N$16330 N$16217 N$16219 "Waveguide Crossing" sch_x=118 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4216 N$16332 N$16334 N$16221 N$16223 "Waveguide Crossing" sch_x=118 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4217 N$16336 N$16338 N$16225 N$16227 "Waveguide Crossing" sch_x=118 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4218 N$16340 N$16342 N$16229 N$16231 "Waveguide Crossing" sch_x=118 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4219 N$16344 N$16346 N$16233 N$16235 "Waveguide Crossing" sch_x=118 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4220 N$16348 N$16350 N$16237 N$16239 "Waveguide Crossing" sch_x=118 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4221 N$16352 N$16354 N$16241 N$16243 "Waveguide Crossing" sch_x=118 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4222 N$16356 N$16358 N$16245 N$16247 "Waveguide Crossing" sch_x=118 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4223 N$16360 N$16362 N$16249 N$16251 "Waveguide Crossing" sch_x=118 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4224 N$16364 N$16366 N$16253 N$16255 "Waveguide Crossing" sch_x=118 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4225 N$16368 N$16370 N$16257 N$16259 "Waveguide Crossing" sch_x=118 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4226 N$16372 N$16374 N$16261 N$16263 "Waveguide Crossing" sch_x=118 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4227 N$16376 N$16378 N$16265 N$16267 "Waveguide Crossing" sch_x=118 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4228 N$16380 N$16382 N$16269 N$16271 "Waveguide Crossing" sch_x=118 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4229 N$16384 N$16386 N$16273 N$16275 "Waveguide Crossing" sch_x=118 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4230 N$16388 N$17909 N$16277 N$16279 "Waveguide Crossing" sch_x=118 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4231 N$17801 N$16390 N$16281 N$16283 "Waveguide Crossing" sch_x=116 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4232 N$16392 N$16394 N$16285 N$16287 "Waveguide Crossing" sch_x=116 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4233 N$16396 N$16398 N$16289 N$16291 "Waveguide Crossing" sch_x=116 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4234 N$16400 N$16402 N$16293 N$16295 "Waveguide Crossing" sch_x=116 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4235 N$16404 N$16406 N$16297 N$16299 "Waveguide Crossing" sch_x=116 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4236 N$16408 N$16410 N$16301 N$16303 "Waveguide Crossing" sch_x=116 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4237 N$16412 N$16414 N$16305 N$16307 "Waveguide Crossing" sch_x=116 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4238 N$16416 N$16418 N$16309 N$16311 "Waveguide Crossing" sch_x=116 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4239 N$16420 N$16422 N$16313 N$16315 "Waveguide Crossing" sch_x=116 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4240 N$16424 N$16426 N$16317 N$16319 "Waveguide Crossing" sch_x=116 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4241 N$16428 N$16430 N$16321 N$16323 "Waveguide Crossing" sch_x=116 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4242 N$16432 N$16434 N$16325 N$16327 "Waveguide Crossing" sch_x=116 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4243 N$16436 N$16438 N$16329 N$16331 "Waveguide Crossing" sch_x=116 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4244 N$16440 N$16442 N$16333 N$16335 "Waveguide Crossing" sch_x=116 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4245 N$16444 N$16446 N$16337 N$16339 "Waveguide Crossing" sch_x=116 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4246 N$16448 N$16450 N$16341 N$16343 "Waveguide Crossing" sch_x=116 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4247 N$16452 N$16454 N$16345 N$16347 "Waveguide Crossing" sch_x=116 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4248 N$16456 N$16458 N$16349 N$16351 "Waveguide Crossing" sch_x=116 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4249 N$16460 N$16462 N$16353 N$16355 "Waveguide Crossing" sch_x=116 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4250 N$16464 N$16466 N$16357 N$16359 "Waveguide Crossing" sch_x=116 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4251 N$16468 N$16470 N$16361 N$16363 "Waveguide Crossing" sch_x=116 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4252 N$16472 N$16474 N$16365 N$16367 "Waveguide Crossing" sch_x=116 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4253 N$16476 N$16478 N$16369 N$16371 "Waveguide Crossing" sch_x=116 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4254 N$16480 N$16482 N$16373 N$16375 "Waveguide Crossing" sch_x=116 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4255 N$16484 N$16486 N$16377 N$16379 "Waveguide Crossing" sch_x=116 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4256 N$16488 N$16490 N$16381 N$16383 "Waveguide Crossing" sch_x=116 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4257 N$16492 N$17907 N$16385 N$16387 "Waveguide Crossing" sch_x=116 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4258 N$17803 N$16494 N$16389 N$16391 "Waveguide Crossing" sch_x=114 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4259 N$16496 N$16498 N$16393 N$16395 "Waveguide Crossing" sch_x=114 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4260 N$16500 N$16502 N$16397 N$16399 "Waveguide Crossing" sch_x=114 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4261 N$16504 N$16506 N$16401 N$16403 "Waveguide Crossing" sch_x=114 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4262 N$16508 N$16510 N$16405 N$16407 "Waveguide Crossing" sch_x=114 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4263 N$16512 N$16514 N$16409 N$16411 "Waveguide Crossing" sch_x=114 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4264 N$16516 N$16518 N$16413 N$16415 "Waveguide Crossing" sch_x=114 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4265 N$16520 N$16522 N$16417 N$16419 "Waveguide Crossing" sch_x=114 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4266 N$16524 N$16526 N$16421 N$16423 "Waveguide Crossing" sch_x=114 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4267 N$16528 N$16530 N$16425 N$16427 "Waveguide Crossing" sch_x=114 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4268 N$16532 N$16534 N$16429 N$16431 "Waveguide Crossing" sch_x=114 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4269 N$16536 N$16538 N$16433 N$16435 "Waveguide Crossing" sch_x=114 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4270 N$16540 N$16542 N$16437 N$16439 "Waveguide Crossing" sch_x=114 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4271 N$16544 N$16546 N$16441 N$16443 "Waveguide Crossing" sch_x=114 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4272 N$16548 N$16550 N$16445 N$16447 "Waveguide Crossing" sch_x=114 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4273 N$16552 N$16554 N$16449 N$16451 "Waveguide Crossing" sch_x=114 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4274 N$16556 N$16558 N$16453 N$16455 "Waveguide Crossing" sch_x=114 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4275 N$16560 N$16562 N$16457 N$16459 "Waveguide Crossing" sch_x=114 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4276 N$16564 N$16566 N$16461 N$16463 "Waveguide Crossing" sch_x=114 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4277 N$16568 N$16570 N$16465 N$16467 "Waveguide Crossing" sch_x=114 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4278 N$16572 N$16574 N$16469 N$16471 "Waveguide Crossing" sch_x=114 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4279 N$16576 N$16578 N$16473 N$16475 "Waveguide Crossing" sch_x=114 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4280 N$16580 N$16582 N$16477 N$16479 "Waveguide Crossing" sch_x=114 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4281 N$16584 N$16586 N$16481 N$16483 "Waveguide Crossing" sch_x=114 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4282 N$16588 N$16590 N$16485 N$16487 "Waveguide Crossing" sch_x=114 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4283 N$16592 N$17905 N$16489 N$16491 "Waveguide Crossing" sch_x=114 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4284 N$17805 N$16594 N$16493 N$16495 "Waveguide Crossing" sch_x=112 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4285 N$16596 N$16598 N$16497 N$16499 "Waveguide Crossing" sch_x=112 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4286 N$16600 N$16602 N$16501 N$16503 "Waveguide Crossing" sch_x=112 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4287 N$16604 N$16606 N$16505 N$16507 "Waveguide Crossing" sch_x=112 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4288 N$16608 N$16610 N$16509 N$16511 "Waveguide Crossing" sch_x=112 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4289 N$16612 N$16614 N$16513 N$16515 "Waveguide Crossing" sch_x=112 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4290 N$16616 N$16618 N$16517 N$16519 "Waveguide Crossing" sch_x=112 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4291 N$16620 N$16622 N$16521 N$16523 "Waveguide Crossing" sch_x=112 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4292 N$16624 N$16626 N$16525 N$16527 "Waveguide Crossing" sch_x=112 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4293 N$16628 N$16630 N$16529 N$16531 "Waveguide Crossing" sch_x=112 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4294 N$16632 N$16634 N$16533 N$16535 "Waveguide Crossing" sch_x=112 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4295 N$16636 N$16638 N$16537 N$16539 "Waveguide Crossing" sch_x=112 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4296 N$16640 N$16642 N$16541 N$16543 "Waveguide Crossing" sch_x=112 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4297 N$16644 N$16646 N$16545 N$16547 "Waveguide Crossing" sch_x=112 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4298 N$16648 N$16650 N$16549 N$16551 "Waveguide Crossing" sch_x=112 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4299 N$16652 N$16654 N$16553 N$16555 "Waveguide Crossing" sch_x=112 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4300 N$16656 N$16658 N$16557 N$16559 "Waveguide Crossing" sch_x=112 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4301 N$16660 N$16662 N$16561 N$16563 "Waveguide Crossing" sch_x=112 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4302 N$16664 N$16666 N$16565 N$16567 "Waveguide Crossing" sch_x=112 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4303 N$16668 N$16670 N$16569 N$16571 "Waveguide Crossing" sch_x=112 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4304 N$16672 N$16674 N$16573 N$16575 "Waveguide Crossing" sch_x=112 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4305 N$16676 N$16678 N$16577 N$16579 "Waveguide Crossing" sch_x=112 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4306 N$16680 N$16682 N$16581 N$16583 "Waveguide Crossing" sch_x=112 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4307 N$16684 N$16686 N$16585 N$16587 "Waveguide Crossing" sch_x=112 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4308 N$16688 N$17903 N$16589 N$16591 "Waveguide Crossing" sch_x=112 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4309 N$17807 N$16690 N$16593 N$16595 "Waveguide Crossing" sch_x=110 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4310 N$16692 N$16694 N$16597 N$16599 "Waveguide Crossing" sch_x=110 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4311 N$16696 N$16698 N$16601 N$16603 "Waveguide Crossing" sch_x=110 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4312 N$16700 N$16702 N$16605 N$16607 "Waveguide Crossing" sch_x=110 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4313 N$16704 N$16706 N$16609 N$16611 "Waveguide Crossing" sch_x=110 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4314 N$16708 N$16710 N$16613 N$16615 "Waveguide Crossing" sch_x=110 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4315 N$16712 N$16714 N$16617 N$16619 "Waveguide Crossing" sch_x=110 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4316 N$16716 N$16718 N$16621 N$16623 "Waveguide Crossing" sch_x=110 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4317 N$16720 N$16722 N$16625 N$16627 "Waveguide Crossing" sch_x=110 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4318 N$16724 N$16726 N$16629 N$16631 "Waveguide Crossing" sch_x=110 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4319 N$16728 N$16730 N$16633 N$16635 "Waveguide Crossing" sch_x=110 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4320 N$16732 N$16734 N$16637 N$16639 "Waveguide Crossing" sch_x=110 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4321 N$16736 N$16738 N$16641 N$16643 "Waveguide Crossing" sch_x=110 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4322 N$16740 N$16742 N$16645 N$16647 "Waveguide Crossing" sch_x=110 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4323 N$16744 N$16746 N$16649 N$16651 "Waveguide Crossing" sch_x=110 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4324 N$16748 N$16750 N$16653 N$16655 "Waveguide Crossing" sch_x=110 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4325 N$16752 N$16754 N$16657 N$16659 "Waveguide Crossing" sch_x=110 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4326 N$16756 N$16758 N$16661 N$16663 "Waveguide Crossing" sch_x=110 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4327 N$16760 N$16762 N$16665 N$16667 "Waveguide Crossing" sch_x=110 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4328 N$16764 N$16766 N$16669 N$16671 "Waveguide Crossing" sch_x=110 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4329 N$16768 N$16770 N$16673 N$16675 "Waveguide Crossing" sch_x=110 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4330 N$16772 N$16774 N$16677 N$16679 "Waveguide Crossing" sch_x=110 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4331 N$16776 N$16778 N$16681 N$16683 "Waveguide Crossing" sch_x=110 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4332 N$16780 N$17901 N$16685 N$16687 "Waveguide Crossing" sch_x=110 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4333 N$17809 N$16782 N$16689 N$16691 "Waveguide Crossing" sch_x=108 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4334 N$16784 N$16786 N$16693 N$16695 "Waveguide Crossing" sch_x=108 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4335 N$16788 N$16790 N$16697 N$16699 "Waveguide Crossing" sch_x=108 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4336 N$16792 N$16794 N$16701 N$16703 "Waveguide Crossing" sch_x=108 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4337 N$16796 N$16798 N$16705 N$16707 "Waveguide Crossing" sch_x=108 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4338 N$16800 N$16802 N$16709 N$16711 "Waveguide Crossing" sch_x=108 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4339 N$16804 N$16806 N$16713 N$16715 "Waveguide Crossing" sch_x=108 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4340 N$16808 N$16810 N$16717 N$16719 "Waveguide Crossing" sch_x=108 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4341 N$16812 N$16814 N$16721 N$16723 "Waveguide Crossing" sch_x=108 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4342 N$16816 N$16818 N$16725 N$16727 "Waveguide Crossing" sch_x=108 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4343 N$16820 N$16822 N$16729 N$16731 "Waveguide Crossing" sch_x=108 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4344 N$16824 N$16826 N$16733 N$16735 "Waveguide Crossing" sch_x=108 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4345 N$16828 N$16830 N$16737 N$16739 "Waveguide Crossing" sch_x=108 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4346 N$16832 N$16834 N$16741 N$16743 "Waveguide Crossing" sch_x=108 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4347 N$16836 N$16838 N$16745 N$16747 "Waveguide Crossing" sch_x=108 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4348 N$16840 N$16842 N$16749 N$16751 "Waveguide Crossing" sch_x=108 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4349 N$16844 N$16846 N$16753 N$16755 "Waveguide Crossing" sch_x=108 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4350 N$16848 N$16850 N$16757 N$16759 "Waveguide Crossing" sch_x=108 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4351 N$16852 N$16854 N$16761 N$16763 "Waveguide Crossing" sch_x=108 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4352 N$16856 N$16858 N$16765 N$16767 "Waveguide Crossing" sch_x=108 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4353 N$16860 N$16862 N$16769 N$16771 "Waveguide Crossing" sch_x=108 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4354 N$16864 N$16866 N$16773 N$16775 "Waveguide Crossing" sch_x=108 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4355 N$16868 N$17899 N$16777 N$16779 "Waveguide Crossing" sch_x=108 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4356 N$17811 N$16870 N$16781 N$16783 "Waveguide Crossing" sch_x=106 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4357 N$16872 N$16874 N$16785 N$16787 "Waveguide Crossing" sch_x=106 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4358 N$16876 N$16878 N$16789 N$16791 "Waveguide Crossing" sch_x=106 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4359 N$16880 N$16882 N$16793 N$16795 "Waveguide Crossing" sch_x=106 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4360 N$16884 N$16886 N$16797 N$16799 "Waveguide Crossing" sch_x=106 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4361 N$16888 N$16890 N$16801 N$16803 "Waveguide Crossing" sch_x=106 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4362 N$16892 N$16894 N$16805 N$16807 "Waveguide Crossing" sch_x=106 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4363 N$16896 N$16898 N$16809 N$16811 "Waveguide Crossing" sch_x=106 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4364 N$16900 N$16902 N$16813 N$16815 "Waveguide Crossing" sch_x=106 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4365 N$16904 N$16906 N$16817 N$16819 "Waveguide Crossing" sch_x=106 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4366 N$16908 N$16910 N$16821 N$16823 "Waveguide Crossing" sch_x=106 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4367 N$16912 N$16914 N$16825 N$16827 "Waveguide Crossing" sch_x=106 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4368 N$16916 N$16918 N$16829 N$16831 "Waveguide Crossing" sch_x=106 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4369 N$16920 N$16922 N$16833 N$16835 "Waveguide Crossing" sch_x=106 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4370 N$16924 N$16926 N$16837 N$16839 "Waveguide Crossing" sch_x=106 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4371 N$16928 N$16930 N$16841 N$16843 "Waveguide Crossing" sch_x=106 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4372 N$16932 N$16934 N$16845 N$16847 "Waveguide Crossing" sch_x=106 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4373 N$16936 N$16938 N$16849 N$16851 "Waveguide Crossing" sch_x=106 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4374 N$16940 N$16942 N$16853 N$16855 "Waveguide Crossing" sch_x=106 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4375 N$16944 N$16946 N$16857 N$16859 "Waveguide Crossing" sch_x=106 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4376 N$16948 N$16950 N$16861 N$16863 "Waveguide Crossing" sch_x=106 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4377 N$16952 N$17897 N$16865 N$16867 "Waveguide Crossing" sch_x=106 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4378 N$17813 N$16954 N$16869 N$16871 "Waveguide Crossing" sch_x=104 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4379 N$16956 N$16958 N$16873 N$16875 "Waveguide Crossing" sch_x=104 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4380 N$16960 N$16962 N$16877 N$16879 "Waveguide Crossing" sch_x=104 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4381 N$16964 N$16966 N$16881 N$16883 "Waveguide Crossing" sch_x=104 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4382 N$16968 N$16970 N$16885 N$16887 "Waveguide Crossing" sch_x=104 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4383 N$16972 N$16974 N$16889 N$16891 "Waveguide Crossing" sch_x=104 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4384 N$16976 N$16978 N$16893 N$16895 "Waveguide Crossing" sch_x=104 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4385 N$16980 N$16982 N$16897 N$16899 "Waveguide Crossing" sch_x=104 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4386 N$16984 N$16986 N$16901 N$16903 "Waveguide Crossing" sch_x=104 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4387 N$16988 N$16990 N$16905 N$16907 "Waveguide Crossing" sch_x=104 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4388 N$16992 N$16994 N$16909 N$16911 "Waveguide Crossing" sch_x=104 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4389 N$16996 N$16998 N$16913 N$16915 "Waveguide Crossing" sch_x=104 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4390 N$17000 N$17002 N$16917 N$16919 "Waveguide Crossing" sch_x=104 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4391 N$17004 N$17006 N$16921 N$16923 "Waveguide Crossing" sch_x=104 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4392 N$17008 N$17010 N$16925 N$16927 "Waveguide Crossing" sch_x=104 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4393 N$17012 N$17014 N$16929 N$16931 "Waveguide Crossing" sch_x=104 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4394 N$17016 N$17018 N$16933 N$16935 "Waveguide Crossing" sch_x=104 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4395 N$17020 N$17022 N$16937 N$16939 "Waveguide Crossing" sch_x=104 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4396 N$17024 N$17026 N$16941 N$16943 "Waveguide Crossing" sch_x=104 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4397 N$17028 N$17030 N$16945 N$16947 "Waveguide Crossing" sch_x=104 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4398 N$17032 N$17895 N$16949 N$16951 "Waveguide Crossing" sch_x=104 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4399 N$17815 N$17034 N$16953 N$16955 "Waveguide Crossing" sch_x=102 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4400 N$17036 N$17038 N$16957 N$16959 "Waveguide Crossing" sch_x=102 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4401 N$17040 N$17042 N$16961 N$16963 "Waveguide Crossing" sch_x=102 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4402 N$17044 N$17046 N$16965 N$16967 "Waveguide Crossing" sch_x=102 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4403 N$17048 N$17050 N$16969 N$16971 "Waveguide Crossing" sch_x=102 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4404 N$17052 N$17054 N$16973 N$16975 "Waveguide Crossing" sch_x=102 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4405 N$17056 N$17058 N$16977 N$16979 "Waveguide Crossing" sch_x=102 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4406 N$17060 N$17062 N$16981 N$16983 "Waveguide Crossing" sch_x=102 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4407 N$17064 N$17066 N$16985 N$16987 "Waveguide Crossing" sch_x=102 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4408 N$17068 N$17070 N$16989 N$16991 "Waveguide Crossing" sch_x=102 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4409 N$17072 N$17074 N$16993 N$16995 "Waveguide Crossing" sch_x=102 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4410 N$17076 N$17078 N$16997 N$16999 "Waveguide Crossing" sch_x=102 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4411 N$17080 N$17082 N$17001 N$17003 "Waveguide Crossing" sch_x=102 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4412 N$17084 N$17086 N$17005 N$17007 "Waveguide Crossing" sch_x=102 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4413 N$17088 N$17090 N$17009 N$17011 "Waveguide Crossing" sch_x=102 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4414 N$17092 N$17094 N$17013 N$17015 "Waveguide Crossing" sch_x=102 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4415 N$17096 N$17098 N$17017 N$17019 "Waveguide Crossing" sch_x=102 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4416 N$17100 N$17102 N$17021 N$17023 "Waveguide Crossing" sch_x=102 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4417 N$17104 N$17106 N$17025 N$17027 "Waveguide Crossing" sch_x=102 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4418 N$17108 N$17893 N$17029 N$17031 "Waveguide Crossing" sch_x=102 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4419 N$17817 N$17110 N$17033 N$17035 "Waveguide Crossing" sch_x=100 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4420 N$17112 N$17114 N$17037 N$17039 "Waveguide Crossing" sch_x=100 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4421 N$17116 N$17118 N$17041 N$17043 "Waveguide Crossing" sch_x=100 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4422 N$17120 N$17122 N$17045 N$17047 "Waveguide Crossing" sch_x=100 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4423 N$17124 N$17126 N$17049 N$17051 "Waveguide Crossing" sch_x=100 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4424 N$17128 N$17130 N$17053 N$17055 "Waveguide Crossing" sch_x=100 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4425 N$17132 N$17134 N$17057 N$17059 "Waveguide Crossing" sch_x=100 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4426 N$17136 N$17138 N$17061 N$17063 "Waveguide Crossing" sch_x=100 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4427 N$17140 N$17142 N$17065 N$17067 "Waveguide Crossing" sch_x=100 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4428 N$17144 N$17146 N$17069 N$17071 "Waveguide Crossing" sch_x=100 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4429 N$17148 N$17150 N$17073 N$17075 "Waveguide Crossing" sch_x=100 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4430 N$17152 N$17154 N$17077 N$17079 "Waveguide Crossing" sch_x=100 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4431 N$17156 N$17158 N$17081 N$17083 "Waveguide Crossing" sch_x=100 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4432 N$17160 N$17162 N$17085 N$17087 "Waveguide Crossing" sch_x=100 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4433 N$17164 N$17166 N$17089 N$17091 "Waveguide Crossing" sch_x=100 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4434 N$17168 N$17170 N$17093 N$17095 "Waveguide Crossing" sch_x=100 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4435 N$17172 N$17174 N$17097 N$17099 "Waveguide Crossing" sch_x=100 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4436 N$17176 N$17178 N$17101 N$17103 "Waveguide Crossing" sch_x=100 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4437 N$17180 N$17891 N$17105 N$17107 "Waveguide Crossing" sch_x=100 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4438 N$17819 N$17182 N$17109 N$17111 "Waveguide Crossing" sch_x=98 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4439 N$17184 N$17186 N$17113 N$17115 "Waveguide Crossing" sch_x=98 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4440 N$17188 N$17190 N$17117 N$17119 "Waveguide Crossing" sch_x=98 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4441 N$17192 N$17194 N$17121 N$17123 "Waveguide Crossing" sch_x=98 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4442 N$17196 N$17198 N$17125 N$17127 "Waveguide Crossing" sch_x=98 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4443 N$17200 N$17202 N$17129 N$17131 "Waveguide Crossing" sch_x=98 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4444 N$17204 N$17206 N$17133 N$17135 "Waveguide Crossing" sch_x=98 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4445 N$17208 N$17210 N$17137 N$17139 "Waveguide Crossing" sch_x=98 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4446 N$17212 N$17214 N$17141 N$17143 "Waveguide Crossing" sch_x=98 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4447 N$17216 N$17218 N$17145 N$17147 "Waveguide Crossing" sch_x=98 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4448 N$17220 N$17222 N$17149 N$17151 "Waveguide Crossing" sch_x=98 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4449 N$17224 N$17226 N$17153 N$17155 "Waveguide Crossing" sch_x=98 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4450 N$17228 N$17230 N$17157 N$17159 "Waveguide Crossing" sch_x=98 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4451 N$17232 N$17234 N$17161 N$17163 "Waveguide Crossing" sch_x=98 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4452 N$17236 N$17238 N$17165 N$17167 "Waveguide Crossing" sch_x=98 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4453 N$17240 N$17242 N$17169 N$17171 "Waveguide Crossing" sch_x=98 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4454 N$17244 N$17246 N$17173 N$17175 "Waveguide Crossing" sch_x=98 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4455 N$17248 N$17889 N$17177 N$17179 "Waveguide Crossing" sch_x=98 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4456 N$17821 N$17250 N$17181 N$17183 "Waveguide Crossing" sch_x=96 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4457 N$17252 N$17254 N$17185 N$17187 "Waveguide Crossing" sch_x=96 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4458 N$17256 N$17258 N$17189 N$17191 "Waveguide Crossing" sch_x=96 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4459 N$17260 N$17262 N$17193 N$17195 "Waveguide Crossing" sch_x=96 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4460 N$17264 N$17266 N$17197 N$17199 "Waveguide Crossing" sch_x=96 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4461 N$17268 N$17270 N$17201 N$17203 "Waveguide Crossing" sch_x=96 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4462 N$17272 N$17274 N$17205 N$17207 "Waveguide Crossing" sch_x=96 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4463 N$17276 N$17278 N$17209 N$17211 "Waveguide Crossing" sch_x=96 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4464 N$17280 N$17282 N$17213 N$17215 "Waveguide Crossing" sch_x=96 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4465 N$17284 N$17286 N$17217 N$17219 "Waveguide Crossing" sch_x=96 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4466 N$17288 N$17290 N$17221 N$17223 "Waveguide Crossing" sch_x=96 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4467 N$17292 N$17294 N$17225 N$17227 "Waveguide Crossing" sch_x=96 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4468 N$17296 N$17298 N$17229 N$17231 "Waveguide Crossing" sch_x=96 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4469 N$17300 N$17302 N$17233 N$17235 "Waveguide Crossing" sch_x=96 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4470 N$17304 N$17306 N$17237 N$17239 "Waveguide Crossing" sch_x=96 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4471 N$17308 N$17310 N$17241 N$17243 "Waveguide Crossing" sch_x=96 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4472 N$17312 N$17887 N$17245 N$17247 "Waveguide Crossing" sch_x=96 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4473 N$17823 N$17314 N$17249 N$17251 "Waveguide Crossing" sch_x=94 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4474 N$17316 N$17318 N$17253 N$17255 "Waveguide Crossing" sch_x=94 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4475 N$17320 N$17322 N$17257 N$17259 "Waveguide Crossing" sch_x=94 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4476 N$17324 N$17326 N$17261 N$17263 "Waveguide Crossing" sch_x=94 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4477 N$17328 N$17330 N$17265 N$17267 "Waveguide Crossing" sch_x=94 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4478 N$17332 N$17334 N$17269 N$17271 "Waveguide Crossing" sch_x=94 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4479 N$17336 N$17338 N$17273 N$17275 "Waveguide Crossing" sch_x=94 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4480 N$17340 N$17342 N$17277 N$17279 "Waveguide Crossing" sch_x=94 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4481 N$17344 N$17346 N$17281 N$17283 "Waveguide Crossing" sch_x=94 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4482 N$17348 N$17350 N$17285 N$17287 "Waveguide Crossing" sch_x=94 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4483 N$17352 N$17354 N$17289 N$17291 "Waveguide Crossing" sch_x=94 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4484 N$17356 N$17358 N$17293 N$17295 "Waveguide Crossing" sch_x=94 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4485 N$17360 N$17362 N$17297 N$17299 "Waveguide Crossing" sch_x=94 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4486 N$17364 N$17366 N$17301 N$17303 "Waveguide Crossing" sch_x=94 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4487 N$17368 N$17370 N$17305 N$17307 "Waveguide Crossing" sch_x=94 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4488 N$17372 N$17885 N$17309 N$17311 "Waveguide Crossing" sch_x=94 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4489 N$17825 N$17374 N$17313 N$17315 "Waveguide Crossing" sch_x=92 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4490 N$17376 N$17378 N$17317 N$17319 "Waveguide Crossing" sch_x=92 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4491 N$17380 N$17382 N$17321 N$17323 "Waveguide Crossing" sch_x=92 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4492 N$17384 N$17386 N$17325 N$17327 "Waveguide Crossing" sch_x=92 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4493 N$17388 N$17390 N$17329 N$17331 "Waveguide Crossing" sch_x=92 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4494 N$17392 N$17394 N$17333 N$17335 "Waveguide Crossing" sch_x=92 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4495 N$17396 N$17398 N$17337 N$17339 "Waveguide Crossing" sch_x=92 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4496 N$17400 N$17402 N$17341 N$17343 "Waveguide Crossing" sch_x=92 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4497 N$17404 N$17406 N$17345 N$17347 "Waveguide Crossing" sch_x=92 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4498 N$17408 N$17410 N$17349 N$17351 "Waveguide Crossing" sch_x=92 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4499 N$17412 N$17414 N$17353 N$17355 "Waveguide Crossing" sch_x=92 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4500 N$17416 N$17418 N$17357 N$17359 "Waveguide Crossing" sch_x=92 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4501 N$17420 N$17422 N$17361 N$17363 "Waveguide Crossing" sch_x=92 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4502 N$17424 N$17426 N$17365 N$17367 "Waveguide Crossing" sch_x=92 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4503 N$17428 N$17883 N$17369 N$17371 "Waveguide Crossing" sch_x=92 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4504 N$17827 N$17430 N$17373 N$17375 "Waveguide Crossing" sch_x=90 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4505 N$17432 N$17434 N$17377 N$17379 "Waveguide Crossing" sch_x=90 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4506 N$17436 N$17438 N$17381 N$17383 "Waveguide Crossing" sch_x=90 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4507 N$17440 N$17442 N$17385 N$17387 "Waveguide Crossing" sch_x=90 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4508 N$17444 N$17446 N$17389 N$17391 "Waveguide Crossing" sch_x=90 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4509 N$17448 N$17450 N$17393 N$17395 "Waveguide Crossing" sch_x=90 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4510 N$17452 N$17454 N$17397 N$17399 "Waveguide Crossing" sch_x=90 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4511 N$17456 N$17458 N$17401 N$17403 "Waveguide Crossing" sch_x=90 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4512 N$17460 N$17462 N$17405 N$17407 "Waveguide Crossing" sch_x=90 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4513 N$17464 N$17466 N$17409 N$17411 "Waveguide Crossing" sch_x=90 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4514 N$17468 N$17470 N$17413 N$17415 "Waveguide Crossing" sch_x=90 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4515 N$17472 N$17474 N$17417 N$17419 "Waveguide Crossing" sch_x=90 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4516 N$17476 N$17478 N$17421 N$17423 "Waveguide Crossing" sch_x=90 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4517 N$17480 N$17881 N$17425 N$17427 "Waveguide Crossing" sch_x=90 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4518 N$17829 N$17482 N$17429 N$17431 "Waveguide Crossing" sch_x=88 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4519 N$17484 N$17486 N$17433 N$17435 "Waveguide Crossing" sch_x=88 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4520 N$17488 N$17490 N$17437 N$17439 "Waveguide Crossing" sch_x=88 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4521 N$17492 N$17494 N$17441 N$17443 "Waveguide Crossing" sch_x=88 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4522 N$17496 N$17498 N$17445 N$17447 "Waveguide Crossing" sch_x=88 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4523 N$17500 N$17502 N$17449 N$17451 "Waveguide Crossing" sch_x=88 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4524 N$17504 N$17506 N$17453 N$17455 "Waveguide Crossing" sch_x=88 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4525 N$17508 N$17510 N$17457 N$17459 "Waveguide Crossing" sch_x=88 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4526 N$17512 N$17514 N$17461 N$17463 "Waveguide Crossing" sch_x=88 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4527 N$17516 N$17518 N$17465 N$17467 "Waveguide Crossing" sch_x=88 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4528 N$17520 N$17522 N$17469 N$17471 "Waveguide Crossing" sch_x=88 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4529 N$17524 N$17526 N$17473 N$17475 "Waveguide Crossing" sch_x=88 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4530 N$17528 N$17879 N$17477 N$17479 "Waveguide Crossing" sch_x=88 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4531 N$17831 N$17530 N$17481 N$17483 "Waveguide Crossing" sch_x=86 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4532 N$17532 N$17534 N$17485 N$17487 "Waveguide Crossing" sch_x=86 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4533 N$17536 N$17538 N$17489 N$17491 "Waveguide Crossing" sch_x=86 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4534 N$17540 N$17542 N$17493 N$17495 "Waveguide Crossing" sch_x=86 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4535 N$17544 N$17546 N$17497 N$17499 "Waveguide Crossing" sch_x=86 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4536 N$17548 N$17550 N$17501 N$17503 "Waveguide Crossing" sch_x=86 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4537 N$17552 N$17554 N$17505 N$17507 "Waveguide Crossing" sch_x=86 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4538 N$17556 N$17558 N$17509 N$17511 "Waveguide Crossing" sch_x=86 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4539 N$17560 N$17562 N$17513 N$17515 "Waveguide Crossing" sch_x=86 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4540 N$17564 N$17566 N$17517 N$17519 "Waveguide Crossing" sch_x=86 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4541 N$17568 N$17570 N$17521 N$17523 "Waveguide Crossing" sch_x=86 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4542 N$17572 N$17877 N$17525 N$17527 "Waveguide Crossing" sch_x=86 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4543 N$17833 N$17574 N$17529 N$17531 "Waveguide Crossing" sch_x=84 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4544 N$17576 N$17578 N$17533 N$17535 "Waveguide Crossing" sch_x=84 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4545 N$17580 N$17582 N$17537 N$17539 "Waveguide Crossing" sch_x=84 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4546 N$17584 N$17586 N$17541 N$17543 "Waveguide Crossing" sch_x=84 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4547 N$17588 N$17590 N$17545 N$17547 "Waveguide Crossing" sch_x=84 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4548 N$17592 N$17594 N$17549 N$17551 "Waveguide Crossing" sch_x=84 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4549 N$17596 N$17598 N$17553 N$17555 "Waveguide Crossing" sch_x=84 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4550 N$17600 N$17602 N$17557 N$17559 "Waveguide Crossing" sch_x=84 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4551 N$17604 N$17606 N$17561 N$17563 "Waveguide Crossing" sch_x=84 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4552 N$17608 N$17610 N$17565 N$17567 "Waveguide Crossing" sch_x=84 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4553 N$17612 N$17875 N$17569 N$17571 "Waveguide Crossing" sch_x=84 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4554 N$17835 N$17614 N$17573 N$17575 "Waveguide Crossing" sch_x=82 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4555 N$17616 N$17618 N$17577 N$17579 "Waveguide Crossing" sch_x=82 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4556 N$17620 N$17622 N$17581 N$17583 "Waveguide Crossing" sch_x=82 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4557 N$17624 N$17626 N$17585 N$17587 "Waveguide Crossing" sch_x=82 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4558 N$17628 N$17630 N$17589 N$17591 "Waveguide Crossing" sch_x=82 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4559 N$17632 N$17634 N$17593 N$17595 "Waveguide Crossing" sch_x=82 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4560 N$17636 N$17638 N$17597 N$17599 "Waveguide Crossing" sch_x=82 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4561 N$17640 N$17642 N$17601 N$17603 "Waveguide Crossing" sch_x=82 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4562 N$17644 N$17646 N$17605 N$17607 "Waveguide Crossing" sch_x=82 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4563 N$17648 N$17873 N$17609 N$17611 "Waveguide Crossing" sch_x=82 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4564 N$17837 N$17650 N$17613 N$17615 "Waveguide Crossing" sch_x=80 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4565 N$17652 N$17654 N$17617 N$17619 "Waveguide Crossing" sch_x=80 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4566 N$17656 N$17658 N$17621 N$17623 "Waveguide Crossing" sch_x=80 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4567 N$17660 N$17662 N$17625 N$17627 "Waveguide Crossing" sch_x=80 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4568 N$17664 N$17666 N$17629 N$17631 "Waveguide Crossing" sch_x=80 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4569 N$17668 N$17670 N$17633 N$17635 "Waveguide Crossing" sch_x=80 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4570 N$17672 N$17674 N$17637 N$17639 "Waveguide Crossing" sch_x=80 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4571 N$17676 N$17678 N$17641 N$17643 "Waveguide Crossing" sch_x=80 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4572 N$17680 N$17871 N$17645 N$17647 "Waveguide Crossing" sch_x=80 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4573 N$17839 N$17682 N$17649 N$17651 "Waveguide Crossing" sch_x=78 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4574 N$17684 N$17686 N$17653 N$17655 "Waveguide Crossing" sch_x=78 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4575 N$17688 N$17690 N$17657 N$17659 "Waveguide Crossing" sch_x=78 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4576 N$17692 N$17694 N$17661 N$17663 "Waveguide Crossing" sch_x=78 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4577 N$17696 N$17698 N$17665 N$17667 "Waveguide Crossing" sch_x=78 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4578 N$17700 N$17702 N$17669 N$17671 "Waveguide Crossing" sch_x=78 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4579 N$17704 N$17706 N$17673 N$17675 "Waveguide Crossing" sch_x=78 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4580 N$17708 N$17869 N$17677 N$17679 "Waveguide Crossing" sch_x=78 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4581 N$17841 N$17710 N$17681 N$17683 "Waveguide Crossing" sch_x=76 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4582 N$17712 N$17714 N$17685 N$17687 "Waveguide Crossing" sch_x=76 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4583 N$17716 N$17718 N$17689 N$17691 "Waveguide Crossing" sch_x=76 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4584 N$17720 N$17722 N$17693 N$17695 "Waveguide Crossing" sch_x=76 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4585 N$17724 N$17726 N$17697 N$17699 "Waveguide Crossing" sch_x=76 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4586 N$17728 N$17730 N$17701 N$17703 "Waveguide Crossing" sch_x=76 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4587 N$17732 N$17867 N$17705 N$17707 "Waveguide Crossing" sch_x=76 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4588 N$17843 N$17734 N$17709 N$17711 "Waveguide Crossing" sch_x=74 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4589 N$17736 N$17738 N$17713 N$17715 "Waveguide Crossing" sch_x=74 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4590 N$17740 N$17742 N$17717 N$17719 "Waveguide Crossing" sch_x=74 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4591 N$17744 N$17746 N$17721 N$17723 "Waveguide Crossing" sch_x=74 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4592 N$17748 N$17750 N$17725 N$17727 "Waveguide Crossing" sch_x=74 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4593 N$17752 N$17865 N$17729 N$17731 "Waveguide Crossing" sch_x=74 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4594 N$17845 N$17754 N$17733 N$17735 "Waveguide Crossing" sch_x=72 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4595 N$17756 N$17758 N$17737 N$17739 "Waveguide Crossing" sch_x=72 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4596 N$17760 N$17762 N$17741 N$17743 "Waveguide Crossing" sch_x=72 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4597 N$17764 N$17766 N$17745 N$17747 "Waveguide Crossing" sch_x=72 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4598 N$17768 N$17863 N$17749 N$17751 "Waveguide Crossing" sch_x=72 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4599 N$17847 N$17770 N$17753 N$17755 "Waveguide Crossing" sch_x=70 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4600 N$17772 N$17774 N$17757 N$17759 "Waveguide Crossing" sch_x=70 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4601 N$17776 N$17778 N$17761 N$17763 "Waveguide Crossing" sch_x=70 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4602 N$17780 N$17861 N$17765 N$17767 "Waveguide Crossing" sch_x=70 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4603 N$17849 N$17782 N$17769 N$17771 "Waveguide Crossing" sch_x=68 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4604 N$17784 N$17786 N$17773 N$17775 "Waveguide Crossing" sch_x=68 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4605 N$17788 N$17859 N$17777 N$17779 "Waveguide Crossing" sch_x=68 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4606 N$17851 N$17790 N$17781 N$17783 "Waveguide Crossing" sch_x=66 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4607 N$17792 N$17857 N$17785 N$17787 "Waveguide Crossing" sch_x=66 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C4608 N$17853 N$17855 N$17789 N$17791 "Waveguide Crossing" sch_x=64 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4081 N$17917 N$15810 N$34432 N$34434 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4082 N$15812 N$15814 N$34436 N$34438 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4083 N$15816 N$15818 N$34440 N$34442 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4084 N$15820 N$15822 N$34444 N$34446 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4085 N$15824 N$15826 N$34448 N$34450 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4086 N$15828 N$15830 N$34452 N$34454 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4087 N$15832 N$15834 N$34456 N$34458 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4088 N$15836 N$15838 N$34460 N$34462 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4089 N$15840 N$15842 N$34464 N$34466 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4090 N$15844 N$15846 N$34468 N$34470 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4091 N$15848 N$15850 N$34472 N$34474 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4092 N$15852 N$15854 N$34476 N$34478 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4093 N$15856 N$15858 N$34480 N$34482 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4094 N$15860 N$15862 N$34484 N$34486 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4095 N$15864 N$15866 N$34488 N$34490 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4096 N$15868 N$15870 N$34492 N$34494 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4097 N$15872 N$15874 N$34496 N$34498 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4098 N$15876 N$15878 N$34500 N$34502 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4099 N$15880 N$15882 N$34504 N$34506 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4100 N$15884 N$15886 N$34508 N$34510 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4101 N$15888 N$15890 N$34512 N$34514 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4102 N$15892 N$15894 N$34516 N$34518 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4103 N$15896 N$15898 N$34520 N$34522 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4104 N$15900 N$15902 N$34524 N$34526 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4105 N$15904 N$15906 N$34528 N$34530 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4106 N$15908 N$15910 N$34532 N$34534 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4107 N$15912 N$15914 N$34536 N$34538 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4108 N$15916 N$15918 N$34540 N$34542 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4109 N$15920 N$15922 N$34544 N$34546 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4110 N$15924 N$15926 N$34548 N$34550 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4111 N$15928 N$15930 N$34552 N$34554 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4112 N$15932 N$17919 N$34556 N$34560 BDC_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6753 N$34305 N$26494 N$26241 N$26243 "Waveguide Crossing" sch_x=252 sch_y=62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6754 N$26496 N$26498 N$26245 N$26247 "Waveguide Crossing" sch_x=252 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6755 N$26500 N$26502 N$26249 N$26251 "Waveguide Crossing" sch_x=252 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6756 N$26504 N$26506 N$26253 N$26255 "Waveguide Crossing" sch_x=252 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6757 N$26508 N$26510 N$26257 N$26259 "Waveguide Crossing" sch_x=252 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6758 N$26512 N$26514 N$26261 N$26263 "Waveguide Crossing" sch_x=252 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6759 N$26516 N$26518 N$26265 N$26267 "Waveguide Crossing" sch_x=252 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6760 N$26520 N$26522 N$26269 N$26271 "Waveguide Crossing" sch_x=252 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6761 N$26524 N$26526 N$26273 N$26275 "Waveguide Crossing" sch_x=252 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6762 N$26528 N$26530 N$26277 N$26279 "Waveguide Crossing" sch_x=252 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6763 N$26532 N$26534 N$26281 N$26283 "Waveguide Crossing" sch_x=252 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6764 N$26536 N$26538 N$26285 N$26287 "Waveguide Crossing" sch_x=252 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6765 N$26540 N$26542 N$26289 N$26291 "Waveguide Crossing" sch_x=252 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6766 N$26544 N$26546 N$26293 N$26295 "Waveguide Crossing" sch_x=252 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6767 N$26548 N$26550 N$26297 N$26299 "Waveguide Crossing" sch_x=252 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6768 N$26552 N$26554 N$26301 N$26303 "Waveguide Crossing" sch_x=252 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6769 N$26556 N$26558 N$26305 N$26307 "Waveguide Crossing" sch_x=252 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6770 N$26560 N$26562 N$26309 N$26311 "Waveguide Crossing" sch_x=252 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6771 N$26564 N$26566 N$26313 N$26315 "Waveguide Crossing" sch_x=252 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6772 N$26568 N$26570 N$26317 N$26319 "Waveguide Crossing" sch_x=252 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6773 N$26572 N$26574 N$26321 N$26323 "Waveguide Crossing" sch_x=252 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6774 N$26576 N$26578 N$26325 N$26327 "Waveguide Crossing" sch_x=252 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6775 N$26580 N$26582 N$26329 N$26331 "Waveguide Crossing" sch_x=252 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6776 N$26584 N$26586 N$26333 N$26335 "Waveguide Crossing" sch_x=252 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6777 N$26588 N$26590 N$26337 N$26339 "Waveguide Crossing" sch_x=252 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6778 N$26592 N$26594 N$26341 N$26343 "Waveguide Crossing" sch_x=252 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6779 N$26596 N$26598 N$26345 N$26347 "Waveguide Crossing" sch_x=252 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6780 N$26600 N$26602 N$26349 N$26351 "Waveguide Crossing" sch_x=252 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6781 N$26604 N$26606 N$26353 N$26355 "Waveguide Crossing" sch_x=252 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6782 N$26608 N$26610 N$26357 N$26359 "Waveguide Crossing" sch_x=252 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6783 N$26612 N$26614 N$26361 N$26363 "Waveguide Crossing" sch_x=252 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6784 N$26616 N$26618 N$26365 N$26367 "Waveguide Crossing" sch_x=252 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6785 N$26620 N$26622 N$26369 N$26371 "Waveguide Crossing" sch_x=252 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6786 N$26624 N$26626 N$26373 N$26375 "Waveguide Crossing" sch_x=252 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6787 N$26628 N$26630 N$26377 N$26379 "Waveguide Crossing" sch_x=252 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6788 N$26632 N$26634 N$26381 N$26383 "Waveguide Crossing" sch_x=252 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6789 N$26636 N$26638 N$26385 N$26387 "Waveguide Crossing" sch_x=252 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6790 N$26640 N$26642 N$26389 N$26391 "Waveguide Crossing" sch_x=252 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6791 N$26644 N$26646 N$26393 N$26395 "Waveguide Crossing" sch_x=252 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6792 N$26648 N$26650 N$26397 N$26399 "Waveguide Crossing" sch_x=252 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6793 N$26652 N$26654 N$26401 N$26403 "Waveguide Crossing" sch_x=252 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6794 N$26656 N$26658 N$26405 N$26407 "Waveguide Crossing" sch_x=252 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6795 N$26660 N$26662 N$26409 N$26411 "Waveguide Crossing" sch_x=252 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6796 N$26664 N$26666 N$26413 N$26415 "Waveguide Crossing" sch_x=252 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6797 N$26668 N$26670 N$26417 N$26419 "Waveguide Crossing" sch_x=252 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6798 N$26672 N$26674 N$26421 N$26423 "Waveguide Crossing" sch_x=252 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6799 N$26676 N$26678 N$26425 N$26427 "Waveguide Crossing" sch_x=252 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6800 N$26680 N$26682 N$26429 N$26431 "Waveguide Crossing" sch_x=252 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6801 N$26684 N$26686 N$26433 N$26435 "Waveguide Crossing" sch_x=252 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6802 N$26688 N$26690 N$26437 N$26439 "Waveguide Crossing" sch_x=252 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6803 N$26692 N$26694 N$26441 N$26443 "Waveguide Crossing" sch_x=252 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6804 N$26696 N$26698 N$26445 N$26447 "Waveguide Crossing" sch_x=252 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6805 N$26700 N$26702 N$26449 N$26451 "Waveguide Crossing" sch_x=252 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6806 N$26704 N$26706 N$26453 N$26455 "Waveguide Crossing" sch_x=252 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6807 N$26708 N$26710 N$26457 N$26459 "Waveguide Crossing" sch_x=252 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6808 N$26712 N$26714 N$26461 N$26463 "Waveguide Crossing" sch_x=252 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6809 N$26716 N$26718 N$26465 N$26467 "Waveguide Crossing" sch_x=252 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6810 N$26720 N$26722 N$26469 N$26471 "Waveguide Crossing" sch_x=252 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6811 N$26724 N$26726 N$26473 N$26475 "Waveguide Crossing" sch_x=252 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6812 N$26728 N$26730 N$26477 N$26479 "Waveguide Crossing" sch_x=252 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6813 N$26732 N$26734 N$26481 N$26483 "Waveguide Crossing" sch_x=252 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6814 N$26736 N$26738 N$26485 N$26487 "Waveguide Crossing" sch_x=252 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6815 N$26740 N$34555 N$26489 N$26491 "Waveguide Crossing" sch_x=252 sch_y=-62 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6816 N$34307 N$26742 N$26493 N$26495 "Waveguide Crossing" sch_x=250 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6817 N$26744 N$26746 N$26497 N$26499 "Waveguide Crossing" sch_x=250 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6818 N$26748 N$26750 N$26501 N$26503 "Waveguide Crossing" sch_x=250 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6819 N$26752 N$26754 N$26505 N$26507 "Waveguide Crossing" sch_x=250 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6820 N$26756 N$26758 N$26509 N$26511 "Waveguide Crossing" sch_x=250 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6821 N$26760 N$26762 N$26513 N$26515 "Waveguide Crossing" sch_x=250 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6822 N$26764 N$26766 N$26517 N$26519 "Waveguide Crossing" sch_x=250 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6823 N$26768 N$26770 N$26521 N$26523 "Waveguide Crossing" sch_x=250 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6824 N$26772 N$26774 N$26525 N$26527 "Waveguide Crossing" sch_x=250 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6825 N$26776 N$26778 N$26529 N$26531 "Waveguide Crossing" sch_x=250 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6826 N$26780 N$26782 N$26533 N$26535 "Waveguide Crossing" sch_x=250 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6827 N$26784 N$26786 N$26537 N$26539 "Waveguide Crossing" sch_x=250 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6828 N$26788 N$26790 N$26541 N$26543 "Waveguide Crossing" sch_x=250 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6829 N$26792 N$26794 N$26545 N$26547 "Waveguide Crossing" sch_x=250 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6830 N$26796 N$26798 N$26549 N$26551 "Waveguide Crossing" sch_x=250 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6831 N$26800 N$26802 N$26553 N$26555 "Waveguide Crossing" sch_x=250 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6832 N$26804 N$26806 N$26557 N$26559 "Waveguide Crossing" sch_x=250 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6833 N$26808 N$26810 N$26561 N$26563 "Waveguide Crossing" sch_x=250 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6834 N$26812 N$26814 N$26565 N$26567 "Waveguide Crossing" sch_x=250 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6835 N$26816 N$26818 N$26569 N$26571 "Waveguide Crossing" sch_x=250 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6836 N$26820 N$26822 N$26573 N$26575 "Waveguide Crossing" sch_x=250 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6837 N$26824 N$26826 N$26577 N$26579 "Waveguide Crossing" sch_x=250 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6838 N$26828 N$26830 N$26581 N$26583 "Waveguide Crossing" sch_x=250 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6839 N$26832 N$26834 N$26585 N$26587 "Waveguide Crossing" sch_x=250 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6840 N$26836 N$26838 N$26589 N$26591 "Waveguide Crossing" sch_x=250 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6841 N$26840 N$26842 N$26593 N$26595 "Waveguide Crossing" sch_x=250 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6842 N$26844 N$26846 N$26597 N$26599 "Waveguide Crossing" sch_x=250 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6843 N$26848 N$26850 N$26601 N$26603 "Waveguide Crossing" sch_x=250 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6844 N$26852 N$26854 N$26605 N$26607 "Waveguide Crossing" sch_x=250 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6845 N$26856 N$26858 N$26609 N$26611 "Waveguide Crossing" sch_x=250 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6846 N$26860 N$26862 N$26613 N$26615 "Waveguide Crossing" sch_x=250 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6847 N$26864 N$26866 N$26617 N$26619 "Waveguide Crossing" sch_x=250 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6848 N$26868 N$26870 N$26621 N$26623 "Waveguide Crossing" sch_x=250 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6849 N$26872 N$26874 N$26625 N$26627 "Waveguide Crossing" sch_x=250 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6850 N$26876 N$26878 N$26629 N$26631 "Waveguide Crossing" sch_x=250 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6851 N$26880 N$26882 N$26633 N$26635 "Waveguide Crossing" sch_x=250 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6852 N$26884 N$26886 N$26637 N$26639 "Waveguide Crossing" sch_x=250 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6853 N$26888 N$26890 N$26641 N$26643 "Waveguide Crossing" sch_x=250 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6854 N$26892 N$26894 N$26645 N$26647 "Waveguide Crossing" sch_x=250 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6855 N$26896 N$26898 N$26649 N$26651 "Waveguide Crossing" sch_x=250 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6856 N$26900 N$26902 N$26653 N$26655 "Waveguide Crossing" sch_x=250 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6857 N$26904 N$26906 N$26657 N$26659 "Waveguide Crossing" sch_x=250 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6858 N$26908 N$26910 N$26661 N$26663 "Waveguide Crossing" sch_x=250 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6859 N$26912 N$26914 N$26665 N$26667 "Waveguide Crossing" sch_x=250 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6860 N$26916 N$26918 N$26669 N$26671 "Waveguide Crossing" sch_x=250 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6861 N$26920 N$26922 N$26673 N$26675 "Waveguide Crossing" sch_x=250 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6862 N$26924 N$26926 N$26677 N$26679 "Waveguide Crossing" sch_x=250 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6863 N$26928 N$26930 N$26681 N$26683 "Waveguide Crossing" sch_x=250 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6864 N$26932 N$26934 N$26685 N$26687 "Waveguide Crossing" sch_x=250 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6865 N$26936 N$26938 N$26689 N$26691 "Waveguide Crossing" sch_x=250 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6866 N$26940 N$26942 N$26693 N$26695 "Waveguide Crossing" sch_x=250 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6867 N$26944 N$26946 N$26697 N$26699 "Waveguide Crossing" sch_x=250 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6868 N$26948 N$26950 N$26701 N$26703 "Waveguide Crossing" sch_x=250 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6869 N$26952 N$26954 N$26705 N$26707 "Waveguide Crossing" sch_x=250 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6870 N$26956 N$26958 N$26709 N$26711 "Waveguide Crossing" sch_x=250 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6871 N$26960 N$26962 N$26713 N$26715 "Waveguide Crossing" sch_x=250 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6872 N$26964 N$26966 N$26717 N$26719 "Waveguide Crossing" sch_x=250 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6873 N$26968 N$26970 N$26721 N$26723 "Waveguide Crossing" sch_x=250 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6874 N$26972 N$26974 N$26725 N$26727 "Waveguide Crossing" sch_x=250 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6875 N$26976 N$26978 N$26729 N$26731 "Waveguide Crossing" sch_x=250 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6876 N$26980 N$26982 N$26733 N$26735 "Waveguide Crossing" sch_x=250 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6877 N$26984 N$34553 N$26737 N$26739 "Waveguide Crossing" sch_x=250 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6878 N$34309 N$26986 N$26741 N$26743 "Waveguide Crossing" sch_x=248 sch_y=60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6879 N$26988 N$26990 N$26745 N$26747 "Waveguide Crossing" sch_x=248 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6880 N$26992 N$26994 N$26749 N$26751 "Waveguide Crossing" sch_x=248 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6881 N$26996 N$26998 N$26753 N$26755 "Waveguide Crossing" sch_x=248 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6882 N$27000 N$27002 N$26757 N$26759 "Waveguide Crossing" sch_x=248 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6883 N$27004 N$27006 N$26761 N$26763 "Waveguide Crossing" sch_x=248 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6884 N$27008 N$27010 N$26765 N$26767 "Waveguide Crossing" sch_x=248 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6885 N$27012 N$27014 N$26769 N$26771 "Waveguide Crossing" sch_x=248 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6886 N$27016 N$27018 N$26773 N$26775 "Waveguide Crossing" sch_x=248 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6887 N$27020 N$27022 N$26777 N$26779 "Waveguide Crossing" sch_x=248 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6888 N$27024 N$27026 N$26781 N$26783 "Waveguide Crossing" sch_x=248 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6889 N$27028 N$27030 N$26785 N$26787 "Waveguide Crossing" sch_x=248 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6890 N$27032 N$27034 N$26789 N$26791 "Waveguide Crossing" sch_x=248 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6891 N$27036 N$27038 N$26793 N$26795 "Waveguide Crossing" sch_x=248 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6892 N$27040 N$27042 N$26797 N$26799 "Waveguide Crossing" sch_x=248 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6893 N$27044 N$27046 N$26801 N$26803 "Waveguide Crossing" sch_x=248 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6894 N$27048 N$27050 N$26805 N$26807 "Waveguide Crossing" sch_x=248 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6895 N$27052 N$27054 N$26809 N$26811 "Waveguide Crossing" sch_x=248 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6896 N$27056 N$27058 N$26813 N$26815 "Waveguide Crossing" sch_x=248 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6897 N$27060 N$27062 N$26817 N$26819 "Waveguide Crossing" sch_x=248 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6898 N$27064 N$27066 N$26821 N$26823 "Waveguide Crossing" sch_x=248 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6899 N$27068 N$27070 N$26825 N$26827 "Waveguide Crossing" sch_x=248 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6900 N$27072 N$27074 N$26829 N$26831 "Waveguide Crossing" sch_x=248 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6901 N$27076 N$27078 N$26833 N$26835 "Waveguide Crossing" sch_x=248 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6902 N$27080 N$27082 N$26837 N$26839 "Waveguide Crossing" sch_x=248 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6903 N$27084 N$27086 N$26841 N$26843 "Waveguide Crossing" sch_x=248 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6904 N$27088 N$27090 N$26845 N$26847 "Waveguide Crossing" sch_x=248 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6905 N$27092 N$27094 N$26849 N$26851 "Waveguide Crossing" sch_x=248 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6906 N$27096 N$27098 N$26853 N$26855 "Waveguide Crossing" sch_x=248 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6907 N$27100 N$27102 N$26857 N$26859 "Waveguide Crossing" sch_x=248 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6908 N$27104 N$27106 N$26861 N$26863 "Waveguide Crossing" sch_x=248 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6909 N$27108 N$27110 N$26865 N$26867 "Waveguide Crossing" sch_x=248 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6910 N$27112 N$27114 N$26869 N$26871 "Waveguide Crossing" sch_x=248 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6911 N$27116 N$27118 N$26873 N$26875 "Waveguide Crossing" sch_x=248 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6912 N$27120 N$27122 N$26877 N$26879 "Waveguide Crossing" sch_x=248 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6913 N$27124 N$27126 N$26881 N$26883 "Waveguide Crossing" sch_x=248 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6914 N$27128 N$27130 N$26885 N$26887 "Waveguide Crossing" sch_x=248 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6915 N$27132 N$27134 N$26889 N$26891 "Waveguide Crossing" sch_x=248 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6916 N$27136 N$27138 N$26893 N$26895 "Waveguide Crossing" sch_x=248 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6917 N$27140 N$27142 N$26897 N$26899 "Waveguide Crossing" sch_x=248 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6918 N$27144 N$27146 N$26901 N$26903 "Waveguide Crossing" sch_x=248 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6919 N$27148 N$27150 N$26905 N$26907 "Waveguide Crossing" sch_x=248 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6920 N$27152 N$27154 N$26909 N$26911 "Waveguide Crossing" sch_x=248 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6921 N$27156 N$27158 N$26913 N$26915 "Waveguide Crossing" sch_x=248 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6922 N$27160 N$27162 N$26917 N$26919 "Waveguide Crossing" sch_x=248 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6923 N$27164 N$27166 N$26921 N$26923 "Waveguide Crossing" sch_x=248 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6924 N$27168 N$27170 N$26925 N$26927 "Waveguide Crossing" sch_x=248 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6925 N$27172 N$27174 N$26929 N$26931 "Waveguide Crossing" sch_x=248 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6926 N$27176 N$27178 N$26933 N$26935 "Waveguide Crossing" sch_x=248 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6927 N$27180 N$27182 N$26937 N$26939 "Waveguide Crossing" sch_x=248 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6928 N$27184 N$27186 N$26941 N$26943 "Waveguide Crossing" sch_x=248 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6929 N$27188 N$27190 N$26945 N$26947 "Waveguide Crossing" sch_x=248 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6930 N$27192 N$27194 N$26949 N$26951 "Waveguide Crossing" sch_x=248 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6931 N$27196 N$27198 N$26953 N$26955 "Waveguide Crossing" sch_x=248 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6932 N$27200 N$27202 N$26957 N$26959 "Waveguide Crossing" sch_x=248 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6933 N$27204 N$27206 N$26961 N$26963 "Waveguide Crossing" sch_x=248 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6934 N$27208 N$27210 N$26965 N$26967 "Waveguide Crossing" sch_x=248 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6935 N$27212 N$27214 N$26969 N$26971 "Waveguide Crossing" sch_x=248 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6936 N$27216 N$27218 N$26973 N$26975 "Waveguide Crossing" sch_x=248 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6937 N$27220 N$27222 N$26977 N$26979 "Waveguide Crossing" sch_x=248 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6938 N$27224 N$34551 N$26981 N$26983 "Waveguide Crossing" sch_x=248 sch_y=-60 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6939 N$34311 N$27226 N$26985 N$26987 "Waveguide Crossing" sch_x=246 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6940 N$27228 N$27230 N$26989 N$26991 "Waveguide Crossing" sch_x=246 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6941 N$27232 N$27234 N$26993 N$26995 "Waveguide Crossing" sch_x=246 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6942 N$27236 N$27238 N$26997 N$26999 "Waveguide Crossing" sch_x=246 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6943 N$27240 N$27242 N$27001 N$27003 "Waveguide Crossing" sch_x=246 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6944 N$27244 N$27246 N$27005 N$27007 "Waveguide Crossing" sch_x=246 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6945 N$27248 N$27250 N$27009 N$27011 "Waveguide Crossing" sch_x=246 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6946 N$27252 N$27254 N$27013 N$27015 "Waveguide Crossing" sch_x=246 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6947 N$27256 N$27258 N$27017 N$27019 "Waveguide Crossing" sch_x=246 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6948 N$27260 N$27262 N$27021 N$27023 "Waveguide Crossing" sch_x=246 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6949 N$27264 N$27266 N$27025 N$27027 "Waveguide Crossing" sch_x=246 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6950 N$27268 N$27270 N$27029 N$27031 "Waveguide Crossing" sch_x=246 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6951 N$27272 N$27274 N$27033 N$27035 "Waveguide Crossing" sch_x=246 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6952 N$27276 N$27278 N$27037 N$27039 "Waveguide Crossing" sch_x=246 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6953 N$27280 N$27282 N$27041 N$27043 "Waveguide Crossing" sch_x=246 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6954 N$27284 N$27286 N$27045 N$27047 "Waveguide Crossing" sch_x=246 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6955 N$27288 N$27290 N$27049 N$27051 "Waveguide Crossing" sch_x=246 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6956 N$27292 N$27294 N$27053 N$27055 "Waveguide Crossing" sch_x=246 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6957 N$27296 N$27298 N$27057 N$27059 "Waveguide Crossing" sch_x=246 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6958 N$27300 N$27302 N$27061 N$27063 "Waveguide Crossing" sch_x=246 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6959 N$27304 N$27306 N$27065 N$27067 "Waveguide Crossing" sch_x=246 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6960 N$27308 N$27310 N$27069 N$27071 "Waveguide Crossing" sch_x=246 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6961 N$27312 N$27314 N$27073 N$27075 "Waveguide Crossing" sch_x=246 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6962 N$27316 N$27318 N$27077 N$27079 "Waveguide Crossing" sch_x=246 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6963 N$27320 N$27322 N$27081 N$27083 "Waveguide Crossing" sch_x=246 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6964 N$27324 N$27326 N$27085 N$27087 "Waveguide Crossing" sch_x=246 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6965 N$27328 N$27330 N$27089 N$27091 "Waveguide Crossing" sch_x=246 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6966 N$27332 N$27334 N$27093 N$27095 "Waveguide Crossing" sch_x=246 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6967 N$27336 N$27338 N$27097 N$27099 "Waveguide Crossing" sch_x=246 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6968 N$27340 N$27342 N$27101 N$27103 "Waveguide Crossing" sch_x=246 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6969 N$27344 N$27346 N$27105 N$27107 "Waveguide Crossing" sch_x=246 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6970 N$27348 N$27350 N$27109 N$27111 "Waveguide Crossing" sch_x=246 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6971 N$27352 N$27354 N$27113 N$27115 "Waveguide Crossing" sch_x=246 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6972 N$27356 N$27358 N$27117 N$27119 "Waveguide Crossing" sch_x=246 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6973 N$27360 N$27362 N$27121 N$27123 "Waveguide Crossing" sch_x=246 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6974 N$27364 N$27366 N$27125 N$27127 "Waveguide Crossing" sch_x=246 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6975 N$27368 N$27370 N$27129 N$27131 "Waveguide Crossing" sch_x=246 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6976 N$27372 N$27374 N$27133 N$27135 "Waveguide Crossing" sch_x=246 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6977 N$27376 N$27378 N$27137 N$27139 "Waveguide Crossing" sch_x=246 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6978 N$27380 N$27382 N$27141 N$27143 "Waveguide Crossing" sch_x=246 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6979 N$27384 N$27386 N$27145 N$27147 "Waveguide Crossing" sch_x=246 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6980 N$27388 N$27390 N$27149 N$27151 "Waveguide Crossing" sch_x=246 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6981 N$27392 N$27394 N$27153 N$27155 "Waveguide Crossing" sch_x=246 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6982 N$27396 N$27398 N$27157 N$27159 "Waveguide Crossing" sch_x=246 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6983 N$27400 N$27402 N$27161 N$27163 "Waveguide Crossing" sch_x=246 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6984 N$27404 N$27406 N$27165 N$27167 "Waveguide Crossing" sch_x=246 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6985 N$27408 N$27410 N$27169 N$27171 "Waveguide Crossing" sch_x=246 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6986 N$27412 N$27414 N$27173 N$27175 "Waveguide Crossing" sch_x=246 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6987 N$27416 N$27418 N$27177 N$27179 "Waveguide Crossing" sch_x=246 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6988 N$27420 N$27422 N$27181 N$27183 "Waveguide Crossing" sch_x=246 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6989 N$27424 N$27426 N$27185 N$27187 "Waveguide Crossing" sch_x=246 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6990 N$27428 N$27430 N$27189 N$27191 "Waveguide Crossing" sch_x=246 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6991 N$27432 N$27434 N$27193 N$27195 "Waveguide Crossing" sch_x=246 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6992 N$27436 N$27438 N$27197 N$27199 "Waveguide Crossing" sch_x=246 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6993 N$27440 N$27442 N$27201 N$27203 "Waveguide Crossing" sch_x=246 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6994 N$27444 N$27446 N$27205 N$27207 "Waveguide Crossing" sch_x=246 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6995 N$27448 N$27450 N$27209 N$27211 "Waveguide Crossing" sch_x=246 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6996 N$27452 N$27454 N$27213 N$27215 "Waveguide Crossing" sch_x=246 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6997 N$27456 N$27458 N$27217 N$27219 "Waveguide Crossing" sch_x=246 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6998 N$27460 N$34549 N$27221 N$27223 "Waveguide Crossing" sch_x=246 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C6999 N$34313 N$27462 N$27225 N$27227 "Waveguide Crossing" sch_x=244 sch_y=58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7000 N$27464 N$27466 N$27229 N$27231 "Waveguide Crossing" sch_x=244 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7001 N$27468 N$27470 N$27233 N$27235 "Waveguide Crossing" sch_x=244 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7002 N$27472 N$27474 N$27237 N$27239 "Waveguide Crossing" sch_x=244 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7003 N$27476 N$27478 N$27241 N$27243 "Waveguide Crossing" sch_x=244 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7004 N$27480 N$27482 N$27245 N$27247 "Waveguide Crossing" sch_x=244 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7005 N$27484 N$27486 N$27249 N$27251 "Waveguide Crossing" sch_x=244 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7006 N$27488 N$27490 N$27253 N$27255 "Waveguide Crossing" sch_x=244 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7007 N$27492 N$27494 N$27257 N$27259 "Waveguide Crossing" sch_x=244 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7008 N$27496 N$27498 N$27261 N$27263 "Waveguide Crossing" sch_x=244 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7009 N$27500 N$27502 N$27265 N$27267 "Waveguide Crossing" sch_x=244 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7010 N$27504 N$27506 N$27269 N$27271 "Waveguide Crossing" sch_x=244 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7011 N$27508 N$27510 N$27273 N$27275 "Waveguide Crossing" sch_x=244 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7012 N$27512 N$27514 N$27277 N$27279 "Waveguide Crossing" sch_x=244 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7013 N$27516 N$27518 N$27281 N$27283 "Waveguide Crossing" sch_x=244 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7014 N$27520 N$27522 N$27285 N$27287 "Waveguide Crossing" sch_x=244 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7015 N$27524 N$27526 N$27289 N$27291 "Waveguide Crossing" sch_x=244 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7016 N$27528 N$27530 N$27293 N$27295 "Waveguide Crossing" sch_x=244 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7017 N$27532 N$27534 N$27297 N$27299 "Waveguide Crossing" sch_x=244 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7018 N$27536 N$27538 N$27301 N$27303 "Waveguide Crossing" sch_x=244 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7019 N$27540 N$27542 N$27305 N$27307 "Waveguide Crossing" sch_x=244 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7020 N$27544 N$27546 N$27309 N$27311 "Waveguide Crossing" sch_x=244 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7021 N$27548 N$27550 N$27313 N$27315 "Waveguide Crossing" sch_x=244 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7022 N$27552 N$27554 N$27317 N$27319 "Waveguide Crossing" sch_x=244 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7023 N$27556 N$27558 N$27321 N$27323 "Waveguide Crossing" sch_x=244 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7024 N$27560 N$27562 N$27325 N$27327 "Waveguide Crossing" sch_x=244 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7025 N$27564 N$27566 N$27329 N$27331 "Waveguide Crossing" sch_x=244 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7026 N$27568 N$27570 N$27333 N$27335 "Waveguide Crossing" sch_x=244 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7027 N$27572 N$27574 N$27337 N$27339 "Waveguide Crossing" sch_x=244 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7028 N$27576 N$27578 N$27341 N$27343 "Waveguide Crossing" sch_x=244 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7029 N$27580 N$27582 N$27345 N$27347 "Waveguide Crossing" sch_x=244 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7030 N$27584 N$27586 N$27349 N$27351 "Waveguide Crossing" sch_x=244 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7031 N$27588 N$27590 N$27353 N$27355 "Waveguide Crossing" sch_x=244 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7032 N$27592 N$27594 N$27357 N$27359 "Waveguide Crossing" sch_x=244 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7033 N$27596 N$27598 N$27361 N$27363 "Waveguide Crossing" sch_x=244 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7034 N$27600 N$27602 N$27365 N$27367 "Waveguide Crossing" sch_x=244 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7035 N$27604 N$27606 N$27369 N$27371 "Waveguide Crossing" sch_x=244 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7036 N$27608 N$27610 N$27373 N$27375 "Waveguide Crossing" sch_x=244 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7037 N$27612 N$27614 N$27377 N$27379 "Waveguide Crossing" sch_x=244 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7038 N$27616 N$27618 N$27381 N$27383 "Waveguide Crossing" sch_x=244 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7039 N$27620 N$27622 N$27385 N$27387 "Waveguide Crossing" sch_x=244 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7040 N$27624 N$27626 N$27389 N$27391 "Waveguide Crossing" sch_x=244 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7041 N$27628 N$27630 N$27393 N$27395 "Waveguide Crossing" sch_x=244 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7042 N$27632 N$27634 N$27397 N$27399 "Waveguide Crossing" sch_x=244 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7043 N$27636 N$27638 N$27401 N$27403 "Waveguide Crossing" sch_x=244 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7044 N$27640 N$27642 N$27405 N$27407 "Waveguide Crossing" sch_x=244 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7045 N$27644 N$27646 N$27409 N$27411 "Waveguide Crossing" sch_x=244 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7046 N$27648 N$27650 N$27413 N$27415 "Waveguide Crossing" sch_x=244 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7047 N$27652 N$27654 N$27417 N$27419 "Waveguide Crossing" sch_x=244 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7048 N$27656 N$27658 N$27421 N$27423 "Waveguide Crossing" sch_x=244 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7049 N$27660 N$27662 N$27425 N$27427 "Waveguide Crossing" sch_x=244 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7050 N$27664 N$27666 N$27429 N$27431 "Waveguide Crossing" sch_x=244 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7051 N$27668 N$27670 N$27433 N$27435 "Waveguide Crossing" sch_x=244 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7052 N$27672 N$27674 N$27437 N$27439 "Waveguide Crossing" sch_x=244 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7053 N$27676 N$27678 N$27441 N$27443 "Waveguide Crossing" sch_x=244 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7054 N$27680 N$27682 N$27445 N$27447 "Waveguide Crossing" sch_x=244 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7055 N$27684 N$27686 N$27449 N$27451 "Waveguide Crossing" sch_x=244 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7056 N$27688 N$27690 N$27453 N$27455 "Waveguide Crossing" sch_x=244 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7057 N$27692 N$34547 N$27457 N$27459 "Waveguide Crossing" sch_x=244 sch_y=-58 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7058 N$34315 N$27694 N$27461 N$27463 "Waveguide Crossing" sch_x=242 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7059 N$27696 N$27698 N$27465 N$27467 "Waveguide Crossing" sch_x=242 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7060 N$27700 N$27702 N$27469 N$27471 "Waveguide Crossing" sch_x=242 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7061 N$27704 N$27706 N$27473 N$27475 "Waveguide Crossing" sch_x=242 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7062 N$27708 N$27710 N$27477 N$27479 "Waveguide Crossing" sch_x=242 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7063 N$27712 N$27714 N$27481 N$27483 "Waveguide Crossing" sch_x=242 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7064 N$27716 N$27718 N$27485 N$27487 "Waveguide Crossing" sch_x=242 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7065 N$27720 N$27722 N$27489 N$27491 "Waveguide Crossing" sch_x=242 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7066 N$27724 N$27726 N$27493 N$27495 "Waveguide Crossing" sch_x=242 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7067 N$27728 N$27730 N$27497 N$27499 "Waveguide Crossing" sch_x=242 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7068 N$27732 N$27734 N$27501 N$27503 "Waveguide Crossing" sch_x=242 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7069 N$27736 N$27738 N$27505 N$27507 "Waveguide Crossing" sch_x=242 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7070 N$27740 N$27742 N$27509 N$27511 "Waveguide Crossing" sch_x=242 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7071 N$27744 N$27746 N$27513 N$27515 "Waveguide Crossing" sch_x=242 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7072 N$27748 N$27750 N$27517 N$27519 "Waveguide Crossing" sch_x=242 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7073 N$27752 N$27754 N$27521 N$27523 "Waveguide Crossing" sch_x=242 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7074 N$27756 N$27758 N$27525 N$27527 "Waveguide Crossing" sch_x=242 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7075 N$27760 N$27762 N$27529 N$27531 "Waveguide Crossing" sch_x=242 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7076 N$27764 N$27766 N$27533 N$27535 "Waveguide Crossing" sch_x=242 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7077 N$27768 N$27770 N$27537 N$27539 "Waveguide Crossing" sch_x=242 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7078 N$27772 N$27774 N$27541 N$27543 "Waveguide Crossing" sch_x=242 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7079 N$27776 N$27778 N$27545 N$27547 "Waveguide Crossing" sch_x=242 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7080 N$27780 N$27782 N$27549 N$27551 "Waveguide Crossing" sch_x=242 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7081 N$27784 N$27786 N$27553 N$27555 "Waveguide Crossing" sch_x=242 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7082 N$27788 N$27790 N$27557 N$27559 "Waveguide Crossing" sch_x=242 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7083 N$27792 N$27794 N$27561 N$27563 "Waveguide Crossing" sch_x=242 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7084 N$27796 N$27798 N$27565 N$27567 "Waveguide Crossing" sch_x=242 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7085 N$27800 N$27802 N$27569 N$27571 "Waveguide Crossing" sch_x=242 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7086 N$27804 N$27806 N$27573 N$27575 "Waveguide Crossing" sch_x=242 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7087 N$27808 N$27810 N$27577 N$27579 "Waveguide Crossing" sch_x=242 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7088 N$27812 N$27814 N$27581 N$27583 "Waveguide Crossing" sch_x=242 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7089 N$27816 N$27818 N$27585 N$27587 "Waveguide Crossing" sch_x=242 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7090 N$27820 N$27822 N$27589 N$27591 "Waveguide Crossing" sch_x=242 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7091 N$27824 N$27826 N$27593 N$27595 "Waveguide Crossing" sch_x=242 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7092 N$27828 N$27830 N$27597 N$27599 "Waveguide Crossing" sch_x=242 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7093 N$27832 N$27834 N$27601 N$27603 "Waveguide Crossing" sch_x=242 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7094 N$27836 N$27838 N$27605 N$27607 "Waveguide Crossing" sch_x=242 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7095 N$27840 N$27842 N$27609 N$27611 "Waveguide Crossing" sch_x=242 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7096 N$27844 N$27846 N$27613 N$27615 "Waveguide Crossing" sch_x=242 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7097 N$27848 N$27850 N$27617 N$27619 "Waveguide Crossing" sch_x=242 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7098 N$27852 N$27854 N$27621 N$27623 "Waveguide Crossing" sch_x=242 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7099 N$27856 N$27858 N$27625 N$27627 "Waveguide Crossing" sch_x=242 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7100 N$27860 N$27862 N$27629 N$27631 "Waveguide Crossing" sch_x=242 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7101 N$27864 N$27866 N$27633 N$27635 "Waveguide Crossing" sch_x=242 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7102 N$27868 N$27870 N$27637 N$27639 "Waveguide Crossing" sch_x=242 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7103 N$27872 N$27874 N$27641 N$27643 "Waveguide Crossing" sch_x=242 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7104 N$27876 N$27878 N$27645 N$27647 "Waveguide Crossing" sch_x=242 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7105 N$27880 N$27882 N$27649 N$27651 "Waveguide Crossing" sch_x=242 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7106 N$27884 N$27886 N$27653 N$27655 "Waveguide Crossing" sch_x=242 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7107 N$27888 N$27890 N$27657 N$27659 "Waveguide Crossing" sch_x=242 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7108 N$27892 N$27894 N$27661 N$27663 "Waveguide Crossing" sch_x=242 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7109 N$27896 N$27898 N$27665 N$27667 "Waveguide Crossing" sch_x=242 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7110 N$27900 N$27902 N$27669 N$27671 "Waveguide Crossing" sch_x=242 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7111 N$27904 N$27906 N$27673 N$27675 "Waveguide Crossing" sch_x=242 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7112 N$27908 N$27910 N$27677 N$27679 "Waveguide Crossing" sch_x=242 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7113 N$27912 N$27914 N$27681 N$27683 "Waveguide Crossing" sch_x=242 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7114 N$27916 N$27918 N$27685 N$27687 "Waveguide Crossing" sch_x=242 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7115 N$27920 N$34545 N$27689 N$27691 "Waveguide Crossing" sch_x=242 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7116 N$34317 N$27922 N$27693 N$27695 "Waveguide Crossing" sch_x=240 sch_y=56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7117 N$27924 N$27926 N$27697 N$27699 "Waveguide Crossing" sch_x=240 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7118 N$27928 N$27930 N$27701 N$27703 "Waveguide Crossing" sch_x=240 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7119 N$27932 N$27934 N$27705 N$27707 "Waveguide Crossing" sch_x=240 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7120 N$27936 N$27938 N$27709 N$27711 "Waveguide Crossing" sch_x=240 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7121 N$27940 N$27942 N$27713 N$27715 "Waveguide Crossing" sch_x=240 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7122 N$27944 N$27946 N$27717 N$27719 "Waveguide Crossing" sch_x=240 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7123 N$27948 N$27950 N$27721 N$27723 "Waveguide Crossing" sch_x=240 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7124 N$27952 N$27954 N$27725 N$27727 "Waveguide Crossing" sch_x=240 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7125 N$27956 N$27958 N$27729 N$27731 "Waveguide Crossing" sch_x=240 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7126 N$27960 N$27962 N$27733 N$27735 "Waveguide Crossing" sch_x=240 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7127 N$27964 N$27966 N$27737 N$27739 "Waveguide Crossing" sch_x=240 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7128 N$27968 N$27970 N$27741 N$27743 "Waveguide Crossing" sch_x=240 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7129 N$27972 N$27974 N$27745 N$27747 "Waveguide Crossing" sch_x=240 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7130 N$27976 N$27978 N$27749 N$27751 "Waveguide Crossing" sch_x=240 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7131 N$27980 N$27982 N$27753 N$27755 "Waveguide Crossing" sch_x=240 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7132 N$27984 N$27986 N$27757 N$27759 "Waveguide Crossing" sch_x=240 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7133 N$27988 N$27990 N$27761 N$27763 "Waveguide Crossing" sch_x=240 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7134 N$27992 N$27994 N$27765 N$27767 "Waveguide Crossing" sch_x=240 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7135 N$27996 N$27998 N$27769 N$27771 "Waveguide Crossing" sch_x=240 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7136 N$28000 N$28002 N$27773 N$27775 "Waveguide Crossing" sch_x=240 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7137 N$28004 N$28006 N$27777 N$27779 "Waveguide Crossing" sch_x=240 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7138 N$28008 N$28010 N$27781 N$27783 "Waveguide Crossing" sch_x=240 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7139 N$28012 N$28014 N$27785 N$27787 "Waveguide Crossing" sch_x=240 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7140 N$28016 N$28018 N$27789 N$27791 "Waveguide Crossing" sch_x=240 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7141 N$28020 N$28022 N$27793 N$27795 "Waveguide Crossing" sch_x=240 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7142 N$28024 N$28026 N$27797 N$27799 "Waveguide Crossing" sch_x=240 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7143 N$28028 N$28030 N$27801 N$27803 "Waveguide Crossing" sch_x=240 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7144 N$28032 N$28034 N$27805 N$27807 "Waveguide Crossing" sch_x=240 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7145 N$28036 N$28038 N$27809 N$27811 "Waveguide Crossing" sch_x=240 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7146 N$28040 N$28042 N$27813 N$27815 "Waveguide Crossing" sch_x=240 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7147 N$28044 N$28046 N$27817 N$27819 "Waveguide Crossing" sch_x=240 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7148 N$28048 N$28050 N$27821 N$27823 "Waveguide Crossing" sch_x=240 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7149 N$28052 N$28054 N$27825 N$27827 "Waveguide Crossing" sch_x=240 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7150 N$28056 N$28058 N$27829 N$27831 "Waveguide Crossing" sch_x=240 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7151 N$28060 N$28062 N$27833 N$27835 "Waveguide Crossing" sch_x=240 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7152 N$28064 N$28066 N$27837 N$27839 "Waveguide Crossing" sch_x=240 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7153 N$28068 N$28070 N$27841 N$27843 "Waveguide Crossing" sch_x=240 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7154 N$28072 N$28074 N$27845 N$27847 "Waveguide Crossing" sch_x=240 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7155 N$28076 N$28078 N$27849 N$27851 "Waveguide Crossing" sch_x=240 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7156 N$28080 N$28082 N$27853 N$27855 "Waveguide Crossing" sch_x=240 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7157 N$28084 N$28086 N$27857 N$27859 "Waveguide Crossing" sch_x=240 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7158 N$28088 N$28090 N$27861 N$27863 "Waveguide Crossing" sch_x=240 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7159 N$28092 N$28094 N$27865 N$27867 "Waveguide Crossing" sch_x=240 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7160 N$28096 N$28098 N$27869 N$27871 "Waveguide Crossing" sch_x=240 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7161 N$28100 N$28102 N$27873 N$27875 "Waveguide Crossing" sch_x=240 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7162 N$28104 N$28106 N$27877 N$27879 "Waveguide Crossing" sch_x=240 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7163 N$28108 N$28110 N$27881 N$27883 "Waveguide Crossing" sch_x=240 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7164 N$28112 N$28114 N$27885 N$27887 "Waveguide Crossing" sch_x=240 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7165 N$28116 N$28118 N$27889 N$27891 "Waveguide Crossing" sch_x=240 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7166 N$28120 N$28122 N$27893 N$27895 "Waveguide Crossing" sch_x=240 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7167 N$28124 N$28126 N$27897 N$27899 "Waveguide Crossing" sch_x=240 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7168 N$28128 N$28130 N$27901 N$27903 "Waveguide Crossing" sch_x=240 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7169 N$28132 N$28134 N$27905 N$27907 "Waveguide Crossing" sch_x=240 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7170 N$28136 N$28138 N$27909 N$27911 "Waveguide Crossing" sch_x=240 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7171 N$28140 N$28142 N$27913 N$27915 "Waveguide Crossing" sch_x=240 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7172 N$28144 N$34543 N$27917 N$27919 "Waveguide Crossing" sch_x=240 sch_y=-56 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7173 N$34319 N$28146 N$27921 N$27923 "Waveguide Crossing" sch_x=238 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7174 N$28148 N$28150 N$27925 N$27927 "Waveguide Crossing" sch_x=238 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7175 N$28152 N$28154 N$27929 N$27931 "Waveguide Crossing" sch_x=238 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7176 N$28156 N$28158 N$27933 N$27935 "Waveguide Crossing" sch_x=238 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7177 N$28160 N$28162 N$27937 N$27939 "Waveguide Crossing" sch_x=238 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7178 N$28164 N$28166 N$27941 N$27943 "Waveguide Crossing" sch_x=238 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7179 N$28168 N$28170 N$27945 N$27947 "Waveguide Crossing" sch_x=238 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7180 N$28172 N$28174 N$27949 N$27951 "Waveguide Crossing" sch_x=238 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7181 N$28176 N$28178 N$27953 N$27955 "Waveguide Crossing" sch_x=238 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7182 N$28180 N$28182 N$27957 N$27959 "Waveguide Crossing" sch_x=238 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7183 N$28184 N$28186 N$27961 N$27963 "Waveguide Crossing" sch_x=238 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7184 N$28188 N$28190 N$27965 N$27967 "Waveguide Crossing" sch_x=238 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7185 N$28192 N$28194 N$27969 N$27971 "Waveguide Crossing" sch_x=238 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7186 N$28196 N$28198 N$27973 N$27975 "Waveguide Crossing" sch_x=238 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7187 N$28200 N$28202 N$27977 N$27979 "Waveguide Crossing" sch_x=238 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7188 N$28204 N$28206 N$27981 N$27983 "Waveguide Crossing" sch_x=238 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7189 N$28208 N$28210 N$27985 N$27987 "Waveguide Crossing" sch_x=238 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7190 N$28212 N$28214 N$27989 N$27991 "Waveguide Crossing" sch_x=238 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7191 N$28216 N$28218 N$27993 N$27995 "Waveguide Crossing" sch_x=238 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7192 N$28220 N$28222 N$27997 N$27999 "Waveguide Crossing" sch_x=238 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7193 N$28224 N$28226 N$28001 N$28003 "Waveguide Crossing" sch_x=238 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7194 N$28228 N$28230 N$28005 N$28007 "Waveguide Crossing" sch_x=238 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7195 N$28232 N$28234 N$28009 N$28011 "Waveguide Crossing" sch_x=238 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7196 N$28236 N$28238 N$28013 N$28015 "Waveguide Crossing" sch_x=238 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7197 N$28240 N$28242 N$28017 N$28019 "Waveguide Crossing" sch_x=238 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7198 N$28244 N$28246 N$28021 N$28023 "Waveguide Crossing" sch_x=238 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7199 N$28248 N$28250 N$28025 N$28027 "Waveguide Crossing" sch_x=238 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7200 N$28252 N$28254 N$28029 N$28031 "Waveguide Crossing" sch_x=238 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7201 N$28256 N$28258 N$28033 N$28035 "Waveguide Crossing" sch_x=238 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7202 N$28260 N$28262 N$28037 N$28039 "Waveguide Crossing" sch_x=238 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7203 N$28264 N$28266 N$28041 N$28043 "Waveguide Crossing" sch_x=238 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7204 N$28268 N$28270 N$28045 N$28047 "Waveguide Crossing" sch_x=238 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7205 N$28272 N$28274 N$28049 N$28051 "Waveguide Crossing" sch_x=238 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7206 N$28276 N$28278 N$28053 N$28055 "Waveguide Crossing" sch_x=238 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7207 N$28280 N$28282 N$28057 N$28059 "Waveguide Crossing" sch_x=238 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7208 N$28284 N$28286 N$28061 N$28063 "Waveguide Crossing" sch_x=238 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7209 N$28288 N$28290 N$28065 N$28067 "Waveguide Crossing" sch_x=238 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7210 N$28292 N$28294 N$28069 N$28071 "Waveguide Crossing" sch_x=238 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7211 N$28296 N$28298 N$28073 N$28075 "Waveguide Crossing" sch_x=238 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7212 N$28300 N$28302 N$28077 N$28079 "Waveguide Crossing" sch_x=238 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7213 N$28304 N$28306 N$28081 N$28083 "Waveguide Crossing" sch_x=238 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7214 N$28308 N$28310 N$28085 N$28087 "Waveguide Crossing" sch_x=238 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7215 N$28312 N$28314 N$28089 N$28091 "Waveguide Crossing" sch_x=238 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7216 N$28316 N$28318 N$28093 N$28095 "Waveguide Crossing" sch_x=238 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7217 N$28320 N$28322 N$28097 N$28099 "Waveguide Crossing" sch_x=238 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7218 N$28324 N$28326 N$28101 N$28103 "Waveguide Crossing" sch_x=238 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7219 N$28328 N$28330 N$28105 N$28107 "Waveguide Crossing" sch_x=238 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7220 N$28332 N$28334 N$28109 N$28111 "Waveguide Crossing" sch_x=238 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7221 N$28336 N$28338 N$28113 N$28115 "Waveguide Crossing" sch_x=238 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7222 N$28340 N$28342 N$28117 N$28119 "Waveguide Crossing" sch_x=238 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7223 N$28344 N$28346 N$28121 N$28123 "Waveguide Crossing" sch_x=238 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7224 N$28348 N$28350 N$28125 N$28127 "Waveguide Crossing" sch_x=238 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7225 N$28352 N$28354 N$28129 N$28131 "Waveguide Crossing" sch_x=238 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7226 N$28356 N$28358 N$28133 N$28135 "Waveguide Crossing" sch_x=238 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7227 N$28360 N$28362 N$28137 N$28139 "Waveguide Crossing" sch_x=238 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7228 N$28364 N$34541 N$28141 N$28143 "Waveguide Crossing" sch_x=238 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7229 N$34321 N$28366 N$28145 N$28147 "Waveguide Crossing" sch_x=236 sch_y=54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7230 N$28368 N$28370 N$28149 N$28151 "Waveguide Crossing" sch_x=236 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7231 N$28372 N$28374 N$28153 N$28155 "Waveguide Crossing" sch_x=236 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7232 N$28376 N$28378 N$28157 N$28159 "Waveguide Crossing" sch_x=236 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7233 N$28380 N$28382 N$28161 N$28163 "Waveguide Crossing" sch_x=236 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7234 N$28384 N$28386 N$28165 N$28167 "Waveguide Crossing" sch_x=236 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7235 N$28388 N$28390 N$28169 N$28171 "Waveguide Crossing" sch_x=236 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7236 N$28392 N$28394 N$28173 N$28175 "Waveguide Crossing" sch_x=236 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7237 N$28396 N$28398 N$28177 N$28179 "Waveguide Crossing" sch_x=236 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7238 N$28400 N$28402 N$28181 N$28183 "Waveguide Crossing" sch_x=236 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7239 N$28404 N$28406 N$28185 N$28187 "Waveguide Crossing" sch_x=236 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7240 N$28408 N$28410 N$28189 N$28191 "Waveguide Crossing" sch_x=236 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7241 N$28412 N$28414 N$28193 N$28195 "Waveguide Crossing" sch_x=236 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7242 N$28416 N$28418 N$28197 N$28199 "Waveguide Crossing" sch_x=236 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7243 N$28420 N$28422 N$28201 N$28203 "Waveguide Crossing" sch_x=236 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7244 N$28424 N$28426 N$28205 N$28207 "Waveguide Crossing" sch_x=236 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7245 N$28428 N$28430 N$28209 N$28211 "Waveguide Crossing" sch_x=236 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7246 N$28432 N$28434 N$28213 N$28215 "Waveguide Crossing" sch_x=236 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7247 N$28436 N$28438 N$28217 N$28219 "Waveguide Crossing" sch_x=236 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7248 N$28440 N$28442 N$28221 N$28223 "Waveguide Crossing" sch_x=236 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7249 N$28444 N$28446 N$28225 N$28227 "Waveguide Crossing" sch_x=236 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7250 N$28448 N$28450 N$28229 N$28231 "Waveguide Crossing" sch_x=236 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7251 N$28452 N$28454 N$28233 N$28235 "Waveguide Crossing" sch_x=236 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7252 N$28456 N$28458 N$28237 N$28239 "Waveguide Crossing" sch_x=236 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7253 N$28460 N$28462 N$28241 N$28243 "Waveguide Crossing" sch_x=236 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7254 N$28464 N$28466 N$28245 N$28247 "Waveguide Crossing" sch_x=236 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7255 N$28468 N$28470 N$28249 N$28251 "Waveguide Crossing" sch_x=236 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7256 N$28472 N$28474 N$28253 N$28255 "Waveguide Crossing" sch_x=236 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7257 N$28476 N$28478 N$28257 N$28259 "Waveguide Crossing" sch_x=236 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7258 N$28480 N$28482 N$28261 N$28263 "Waveguide Crossing" sch_x=236 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7259 N$28484 N$28486 N$28265 N$28267 "Waveguide Crossing" sch_x=236 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7260 N$28488 N$28490 N$28269 N$28271 "Waveguide Crossing" sch_x=236 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7261 N$28492 N$28494 N$28273 N$28275 "Waveguide Crossing" sch_x=236 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7262 N$28496 N$28498 N$28277 N$28279 "Waveguide Crossing" sch_x=236 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7263 N$28500 N$28502 N$28281 N$28283 "Waveguide Crossing" sch_x=236 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7264 N$28504 N$28506 N$28285 N$28287 "Waveguide Crossing" sch_x=236 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7265 N$28508 N$28510 N$28289 N$28291 "Waveguide Crossing" sch_x=236 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7266 N$28512 N$28514 N$28293 N$28295 "Waveguide Crossing" sch_x=236 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7267 N$28516 N$28518 N$28297 N$28299 "Waveguide Crossing" sch_x=236 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7268 N$28520 N$28522 N$28301 N$28303 "Waveguide Crossing" sch_x=236 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7269 N$28524 N$28526 N$28305 N$28307 "Waveguide Crossing" sch_x=236 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7270 N$28528 N$28530 N$28309 N$28311 "Waveguide Crossing" sch_x=236 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7271 N$28532 N$28534 N$28313 N$28315 "Waveguide Crossing" sch_x=236 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7272 N$28536 N$28538 N$28317 N$28319 "Waveguide Crossing" sch_x=236 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7273 N$28540 N$28542 N$28321 N$28323 "Waveguide Crossing" sch_x=236 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7274 N$28544 N$28546 N$28325 N$28327 "Waveguide Crossing" sch_x=236 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7275 N$28548 N$28550 N$28329 N$28331 "Waveguide Crossing" sch_x=236 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7276 N$28552 N$28554 N$28333 N$28335 "Waveguide Crossing" sch_x=236 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7277 N$28556 N$28558 N$28337 N$28339 "Waveguide Crossing" sch_x=236 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7278 N$28560 N$28562 N$28341 N$28343 "Waveguide Crossing" sch_x=236 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7279 N$28564 N$28566 N$28345 N$28347 "Waveguide Crossing" sch_x=236 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7280 N$28568 N$28570 N$28349 N$28351 "Waveguide Crossing" sch_x=236 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7281 N$28572 N$28574 N$28353 N$28355 "Waveguide Crossing" sch_x=236 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7282 N$28576 N$28578 N$28357 N$28359 "Waveguide Crossing" sch_x=236 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7283 N$28580 N$34539 N$28361 N$28363 "Waveguide Crossing" sch_x=236 sch_y=-54 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7284 N$34323 N$28582 N$28365 N$28367 "Waveguide Crossing" sch_x=234 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7285 N$28584 N$28586 N$28369 N$28371 "Waveguide Crossing" sch_x=234 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7286 N$28588 N$28590 N$28373 N$28375 "Waveguide Crossing" sch_x=234 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7287 N$28592 N$28594 N$28377 N$28379 "Waveguide Crossing" sch_x=234 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7288 N$28596 N$28598 N$28381 N$28383 "Waveguide Crossing" sch_x=234 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7289 N$28600 N$28602 N$28385 N$28387 "Waveguide Crossing" sch_x=234 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7290 N$28604 N$28606 N$28389 N$28391 "Waveguide Crossing" sch_x=234 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7291 N$28608 N$28610 N$28393 N$28395 "Waveguide Crossing" sch_x=234 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7292 N$28612 N$28614 N$28397 N$28399 "Waveguide Crossing" sch_x=234 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7293 N$28616 N$28618 N$28401 N$28403 "Waveguide Crossing" sch_x=234 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7294 N$28620 N$28622 N$28405 N$28407 "Waveguide Crossing" sch_x=234 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7295 N$28624 N$28626 N$28409 N$28411 "Waveguide Crossing" sch_x=234 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7296 N$28628 N$28630 N$28413 N$28415 "Waveguide Crossing" sch_x=234 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7297 N$28632 N$28634 N$28417 N$28419 "Waveguide Crossing" sch_x=234 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7298 N$28636 N$28638 N$28421 N$28423 "Waveguide Crossing" sch_x=234 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7299 N$28640 N$28642 N$28425 N$28427 "Waveguide Crossing" sch_x=234 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7300 N$28644 N$28646 N$28429 N$28431 "Waveguide Crossing" sch_x=234 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7301 N$28648 N$28650 N$28433 N$28435 "Waveguide Crossing" sch_x=234 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7302 N$28652 N$28654 N$28437 N$28439 "Waveguide Crossing" sch_x=234 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7303 N$28656 N$28658 N$28441 N$28443 "Waveguide Crossing" sch_x=234 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7304 N$28660 N$28662 N$28445 N$28447 "Waveguide Crossing" sch_x=234 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7305 N$28664 N$28666 N$28449 N$28451 "Waveguide Crossing" sch_x=234 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7306 N$28668 N$28670 N$28453 N$28455 "Waveguide Crossing" sch_x=234 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7307 N$28672 N$28674 N$28457 N$28459 "Waveguide Crossing" sch_x=234 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7308 N$28676 N$28678 N$28461 N$28463 "Waveguide Crossing" sch_x=234 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7309 N$28680 N$28682 N$28465 N$28467 "Waveguide Crossing" sch_x=234 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7310 N$28684 N$28686 N$28469 N$28471 "Waveguide Crossing" sch_x=234 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7311 N$28688 N$28690 N$28473 N$28475 "Waveguide Crossing" sch_x=234 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7312 N$28692 N$28694 N$28477 N$28479 "Waveguide Crossing" sch_x=234 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7313 N$28696 N$28698 N$28481 N$28483 "Waveguide Crossing" sch_x=234 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7314 N$28700 N$28702 N$28485 N$28487 "Waveguide Crossing" sch_x=234 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7315 N$28704 N$28706 N$28489 N$28491 "Waveguide Crossing" sch_x=234 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7316 N$28708 N$28710 N$28493 N$28495 "Waveguide Crossing" sch_x=234 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7317 N$28712 N$28714 N$28497 N$28499 "Waveguide Crossing" sch_x=234 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7318 N$28716 N$28718 N$28501 N$28503 "Waveguide Crossing" sch_x=234 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7319 N$28720 N$28722 N$28505 N$28507 "Waveguide Crossing" sch_x=234 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7320 N$28724 N$28726 N$28509 N$28511 "Waveguide Crossing" sch_x=234 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7321 N$28728 N$28730 N$28513 N$28515 "Waveguide Crossing" sch_x=234 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7322 N$28732 N$28734 N$28517 N$28519 "Waveguide Crossing" sch_x=234 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7323 N$28736 N$28738 N$28521 N$28523 "Waveguide Crossing" sch_x=234 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7324 N$28740 N$28742 N$28525 N$28527 "Waveguide Crossing" sch_x=234 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7325 N$28744 N$28746 N$28529 N$28531 "Waveguide Crossing" sch_x=234 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7326 N$28748 N$28750 N$28533 N$28535 "Waveguide Crossing" sch_x=234 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7327 N$28752 N$28754 N$28537 N$28539 "Waveguide Crossing" sch_x=234 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7328 N$28756 N$28758 N$28541 N$28543 "Waveguide Crossing" sch_x=234 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7329 N$28760 N$28762 N$28545 N$28547 "Waveguide Crossing" sch_x=234 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7330 N$28764 N$28766 N$28549 N$28551 "Waveguide Crossing" sch_x=234 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7331 N$28768 N$28770 N$28553 N$28555 "Waveguide Crossing" sch_x=234 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7332 N$28772 N$28774 N$28557 N$28559 "Waveguide Crossing" sch_x=234 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7333 N$28776 N$28778 N$28561 N$28563 "Waveguide Crossing" sch_x=234 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7334 N$28780 N$28782 N$28565 N$28567 "Waveguide Crossing" sch_x=234 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7335 N$28784 N$28786 N$28569 N$28571 "Waveguide Crossing" sch_x=234 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7336 N$28788 N$28790 N$28573 N$28575 "Waveguide Crossing" sch_x=234 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7337 N$28792 N$34537 N$28577 N$28579 "Waveguide Crossing" sch_x=234 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7338 N$34325 N$28794 N$28581 N$28583 "Waveguide Crossing" sch_x=232 sch_y=52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7339 N$28796 N$28798 N$28585 N$28587 "Waveguide Crossing" sch_x=232 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7340 N$28800 N$28802 N$28589 N$28591 "Waveguide Crossing" sch_x=232 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7341 N$28804 N$28806 N$28593 N$28595 "Waveguide Crossing" sch_x=232 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7342 N$28808 N$28810 N$28597 N$28599 "Waveguide Crossing" sch_x=232 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7343 N$28812 N$28814 N$28601 N$28603 "Waveguide Crossing" sch_x=232 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7344 N$28816 N$28818 N$28605 N$28607 "Waveguide Crossing" sch_x=232 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7345 N$28820 N$28822 N$28609 N$28611 "Waveguide Crossing" sch_x=232 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7346 N$28824 N$28826 N$28613 N$28615 "Waveguide Crossing" sch_x=232 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7347 N$28828 N$28830 N$28617 N$28619 "Waveguide Crossing" sch_x=232 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7348 N$28832 N$28834 N$28621 N$28623 "Waveguide Crossing" sch_x=232 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7349 N$28836 N$28838 N$28625 N$28627 "Waveguide Crossing" sch_x=232 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7350 N$28840 N$28842 N$28629 N$28631 "Waveguide Crossing" sch_x=232 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7351 N$28844 N$28846 N$28633 N$28635 "Waveguide Crossing" sch_x=232 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7352 N$28848 N$28850 N$28637 N$28639 "Waveguide Crossing" sch_x=232 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7353 N$28852 N$28854 N$28641 N$28643 "Waveguide Crossing" sch_x=232 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7354 N$28856 N$28858 N$28645 N$28647 "Waveguide Crossing" sch_x=232 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7355 N$28860 N$28862 N$28649 N$28651 "Waveguide Crossing" sch_x=232 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7356 N$28864 N$28866 N$28653 N$28655 "Waveguide Crossing" sch_x=232 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7357 N$28868 N$28870 N$28657 N$28659 "Waveguide Crossing" sch_x=232 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7358 N$28872 N$28874 N$28661 N$28663 "Waveguide Crossing" sch_x=232 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7359 N$28876 N$28878 N$28665 N$28667 "Waveguide Crossing" sch_x=232 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7360 N$28880 N$28882 N$28669 N$28671 "Waveguide Crossing" sch_x=232 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7361 N$28884 N$28886 N$28673 N$28675 "Waveguide Crossing" sch_x=232 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7362 N$28888 N$28890 N$28677 N$28679 "Waveguide Crossing" sch_x=232 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7363 N$28892 N$28894 N$28681 N$28683 "Waveguide Crossing" sch_x=232 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7364 N$28896 N$28898 N$28685 N$28687 "Waveguide Crossing" sch_x=232 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7365 N$28900 N$28902 N$28689 N$28691 "Waveguide Crossing" sch_x=232 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7366 N$28904 N$28906 N$28693 N$28695 "Waveguide Crossing" sch_x=232 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7367 N$28908 N$28910 N$28697 N$28699 "Waveguide Crossing" sch_x=232 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7368 N$28912 N$28914 N$28701 N$28703 "Waveguide Crossing" sch_x=232 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7369 N$28916 N$28918 N$28705 N$28707 "Waveguide Crossing" sch_x=232 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7370 N$28920 N$28922 N$28709 N$28711 "Waveguide Crossing" sch_x=232 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7371 N$28924 N$28926 N$28713 N$28715 "Waveguide Crossing" sch_x=232 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7372 N$28928 N$28930 N$28717 N$28719 "Waveguide Crossing" sch_x=232 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7373 N$28932 N$28934 N$28721 N$28723 "Waveguide Crossing" sch_x=232 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7374 N$28936 N$28938 N$28725 N$28727 "Waveguide Crossing" sch_x=232 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7375 N$28940 N$28942 N$28729 N$28731 "Waveguide Crossing" sch_x=232 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7376 N$28944 N$28946 N$28733 N$28735 "Waveguide Crossing" sch_x=232 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7377 N$28948 N$28950 N$28737 N$28739 "Waveguide Crossing" sch_x=232 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7378 N$28952 N$28954 N$28741 N$28743 "Waveguide Crossing" sch_x=232 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7379 N$28956 N$28958 N$28745 N$28747 "Waveguide Crossing" sch_x=232 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7380 N$28960 N$28962 N$28749 N$28751 "Waveguide Crossing" sch_x=232 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7381 N$28964 N$28966 N$28753 N$28755 "Waveguide Crossing" sch_x=232 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7382 N$28968 N$28970 N$28757 N$28759 "Waveguide Crossing" sch_x=232 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7383 N$28972 N$28974 N$28761 N$28763 "Waveguide Crossing" sch_x=232 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7384 N$28976 N$28978 N$28765 N$28767 "Waveguide Crossing" sch_x=232 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7385 N$28980 N$28982 N$28769 N$28771 "Waveguide Crossing" sch_x=232 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7386 N$28984 N$28986 N$28773 N$28775 "Waveguide Crossing" sch_x=232 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7387 N$28988 N$28990 N$28777 N$28779 "Waveguide Crossing" sch_x=232 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7388 N$28992 N$28994 N$28781 N$28783 "Waveguide Crossing" sch_x=232 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7389 N$28996 N$28998 N$28785 N$28787 "Waveguide Crossing" sch_x=232 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7390 N$29000 N$34535 N$28789 N$28791 "Waveguide Crossing" sch_x=232 sch_y=-52 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7391 N$34327 N$29002 N$28793 N$28795 "Waveguide Crossing" sch_x=230 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7392 N$29004 N$29006 N$28797 N$28799 "Waveguide Crossing" sch_x=230 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7393 N$29008 N$29010 N$28801 N$28803 "Waveguide Crossing" sch_x=230 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7394 N$29012 N$29014 N$28805 N$28807 "Waveguide Crossing" sch_x=230 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7395 N$29016 N$29018 N$28809 N$28811 "Waveguide Crossing" sch_x=230 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7396 N$29020 N$29022 N$28813 N$28815 "Waveguide Crossing" sch_x=230 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7397 N$29024 N$29026 N$28817 N$28819 "Waveguide Crossing" sch_x=230 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7398 N$29028 N$29030 N$28821 N$28823 "Waveguide Crossing" sch_x=230 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7399 N$29032 N$29034 N$28825 N$28827 "Waveguide Crossing" sch_x=230 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7400 N$29036 N$29038 N$28829 N$28831 "Waveguide Crossing" sch_x=230 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7401 N$29040 N$29042 N$28833 N$28835 "Waveguide Crossing" sch_x=230 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7402 N$29044 N$29046 N$28837 N$28839 "Waveguide Crossing" sch_x=230 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7403 N$29048 N$29050 N$28841 N$28843 "Waveguide Crossing" sch_x=230 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7404 N$29052 N$29054 N$28845 N$28847 "Waveguide Crossing" sch_x=230 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7405 N$29056 N$29058 N$28849 N$28851 "Waveguide Crossing" sch_x=230 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7406 N$29060 N$29062 N$28853 N$28855 "Waveguide Crossing" sch_x=230 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7407 N$29064 N$29066 N$28857 N$28859 "Waveguide Crossing" sch_x=230 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7408 N$29068 N$29070 N$28861 N$28863 "Waveguide Crossing" sch_x=230 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7409 N$29072 N$29074 N$28865 N$28867 "Waveguide Crossing" sch_x=230 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7410 N$29076 N$29078 N$28869 N$28871 "Waveguide Crossing" sch_x=230 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7411 N$29080 N$29082 N$28873 N$28875 "Waveguide Crossing" sch_x=230 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7412 N$29084 N$29086 N$28877 N$28879 "Waveguide Crossing" sch_x=230 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7413 N$29088 N$29090 N$28881 N$28883 "Waveguide Crossing" sch_x=230 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7414 N$29092 N$29094 N$28885 N$28887 "Waveguide Crossing" sch_x=230 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7415 N$29096 N$29098 N$28889 N$28891 "Waveguide Crossing" sch_x=230 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7416 N$29100 N$29102 N$28893 N$28895 "Waveguide Crossing" sch_x=230 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7417 N$29104 N$29106 N$28897 N$28899 "Waveguide Crossing" sch_x=230 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7418 N$29108 N$29110 N$28901 N$28903 "Waveguide Crossing" sch_x=230 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7419 N$29112 N$29114 N$28905 N$28907 "Waveguide Crossing" sch_x=230 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7420 N$29116 N$29118 N$28909 N$28911 "Waveguide Crossing" sch_x=230 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7421 N$29120 N$29122 N$28913 N$28915 "Waveguide Crossing" sch_x=230 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7422 N$29124 N$29126 N$28917 N$28919 "Waveguide Crossing" sch_x=230 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7423 N$29128 N$29130 N$28921 N$28923 "Waveguide Crossing" sch_x=230 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7424 N$29132 N$29134 N$28925 N$28927 "Waveguide Crossing" sch_x=230 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7425 N$29136 N$29138 N$28929 N$28931 "Waveguide Crossing" sch_x=230 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7426 N$29140 N$29142 N$28933 N$28935 "Waveguide Crossing" sch_x=230 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7427 N$29144 N$29146 N$28937 N$28939 "Waveguide Crossing" sch_x=230 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7428 N$29148 N$29150 N$28941 N$28943 "Waveguide Crossing" sch_x=230 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7429 N$29152 N$29154 N$28945 N$28947 "Waveguide Crossing" sch_x=230 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7430 N$29156 N$29158 N$28949 N$28951 "Waveguide Crossing" sch_x=230 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7431 N$29160 N$29162 N$28953 N$28955 "Waveguide Crossing" sch_x=230 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7432 N$29164 N$29166 N$28957 N$28959 "Waveguide Crossing" sch_x=230 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7433 N$29168 N$29170 N$28961 N$28963 "Waveguide Crossing" sch_x=230 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7434 N$29172 N$29174 N$28965 N$28967 "Waveguide Crossing" sch_x=230 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7435 N$29176 N$29178 N$28969 N$28971 "Waveguide Crossing" sch_x=230 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7436 N$29180 N$29182 N$28973 N$28975 "Waveguide Crossing" sch_x=230 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7437 N$29184 N$29186 N$28977 N$28979 "Waveguide Crossing" sch_x=230 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7438 N$29188 N$29190 N$28981 N$28983 "Waveguide Crossing" sch_x=230 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7439 N$29192 N$29194 N$28985 N$28987 "Waveguide Crossing" sch_x=230 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7440 N$29196 N$29198 N$28989 N$28991 "Waveguide Crossing" sch_x=230 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7441 N$29200 N$29202 N$28993 N$28995 "Waveguide Crossing" sch_x=230 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7442 N$29204 N$34533 N$28997 N$28999 "Waveguide Crossing" sch_x=230 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7443 N$34329 N$29206 N$29001 N$29003 "Waveguide Crossing" sch_x=228 sch_y=50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7444 N$29208 N$29210 N$29005 N$29007 "Waveguide Crossing" sch_x=228 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7445 N$29212 N$29214 N$29009 N$29011 "Waveguide Crossing" sch_x=228 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7446 N$29216 N$29218 N$29013 N$29015 "Waveguide Crossing" sch_x=228 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7447 N$29220 N$29222 N$29017 N$29019 "Waveguide Crossing" sch_x=228 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7448 N$29224 N$29226 N$29021 N$29023 "Waveguide Crossing" sch_x=228 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7449 N$29228 N$29230 N$29025 N$29027 "Waveguide Crossing" sch_x=228 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7450 N$29232 N$29234 N$29029 N$29031 "Waveguide Crossing" sch_x=228 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7451 N$29236 N$29238 N$29033 N$29035 "Waveguide Crossing" sch_x=228 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7452 N$29240 N$29242 N$29037 N$29039 "Waveguide Crossing" sch_x=228 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7453 N$29244 N$29246 N$29041 N$29043 "Waveguide Crossing" sch_x=228 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7454 N$29248 N$29250 N$29045 N$29047 "Waveguide Crossing" sch_x=228 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7455 N$29252 N$29254 N$29049 N$29051 "Waveguide Crossing" sch_x=228 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7456 N$29256 N$29258 N$29053 N$29055 "Waveguide Crossing" sch_x=228 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7457 N$29260 N$29262 N$29057 N$29059 "Waveguide Crossing" sch_x=228 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7458 N$29264 N$29266 N$29061 N$29063 "Waveguide Crossing" sch_x=228 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7459 N$29268 N$29270 N$29065 N$29067 "Waveguide Crossing" sch_x=228 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7460 N$29272 N$29274 N$29069 N$29071 "Waveguide Crossing" sch_x=228 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7461 N$29276 N$29278 N$29073 N$29075 "Waveguide Crossing" sch_x=228 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7462 N$29280 N$29282 N$29077 N$29079 "Waveguide Crossing" sch_x=228 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7463 N$29284 N$29286 N$29081 N$29083 "Waveguide Crossing" sch_x=228 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7464 N$29288 N$29290 N$29085 N$29087 "Waveguide Crossing" sch_x=228 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7465 N$29292 N$29294 N$29089 N$29091 "Waveguide Crossing" sch_x=228 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7466 N$29296 N$29298 N$29093 N$29095 "Waveguide Crossing" sch_x=228 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7467 N$29300 N$29302 N$29097 N$29099 "Waveguide Crossing" sch_x=228 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7468 N$29304 N$29306 N$29101 N$29103 "Waveguide Crossing" sch_x=228 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7469 N$29308 N$29310 N$29105 N$29107 "Waveguide Crossing" sch_x=228 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7470 N$29312 N$29314 N$29109 N$29111 "Waveguide Crossing" sch_x=228 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7471 N$29316 N$29318 N$29113 N$29115 "Waveguide Crossing" sch_x=228 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7472 N$29320 N$29322 N$29117 N$29119 "Waveguide Crossing" sch_x=228 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7473 N$29324 N$29326 N$29121 N$29123 "Waveguide Crossing" sch_x=228 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7474 N$29328 N$29330 N$29125 N$29127 "Waveguide Crossing" sch_x=228 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7475 N$29332 N$29334 N$29129 N$29131 "Waveguide Crossing" sch_x=228 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7476 N$29336 N$29338 N$29133 N$29135 "Waveguide Crossing" sch_x=228 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7477 N$29340 N$29342 N$29137 N$29139 "Waveguide Crossing" sch_x=228 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7478 N$29344 N$29346 N$29141 N$29143 "Waveguide Crossing" sch_x=228 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7479 N$29348 N$29350 N$29145 N$29147 "Waveguide Crossing" sch_x=228 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7480 N$29352 N$29354 N$29149 N$29151 "Waveguide Crossing" sch_x=228 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7481 N$29356 N$29358 N$29153 N$29155 "Waveguide Crossing" sch_x=228 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7482 N$29360 N$29362 N$29157 N$29159 "Waveguide Crossing" sch_x=228 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7483 N$29364 N$29366 N$29161 N$29163 "Waveguide Crossing" sch_x=228 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7484 N$29368 N$29370 N$29165 N$29167 "Waveguide Crossing" sch_x=228 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7485 N$29372 N$29374 N$29169 N$29171 "Waveguide Crossing" sch_x=228 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7486 N$29376 N$29378 N$29173 N$29175 "Waveguide Crossing" sch_x=228 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7487 N$29380 N$29382 N$29177 N$29179 "Waveguide Crossing" sch_x=228 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7488 N$29384 N$29386 N$29181 N$29183 "Waveguide Crossing" sch_x=228 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7489 N$29388 N$29390 N$29185 N$29187 "Waveguide Crossing" sch_x=228 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7490 N$29392 N$29394 N$29189 N$29191 "Waveguide Crossing" sch_x=228 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7491 N$29396 N$29398 N$29193 N$29195 "Waveguide Crossing" sch_x=228 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7492 N$29400 N$29402 N$29197 N$29199 "Waveguide Crossing" sch_x=228 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7493 N$29404 N$34531 N$29201 N$29203 "Waveguide Crossing" sch_x=228 sch_y=-50 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7494 N$34331 N$29406 N$29205 N$29207 "Waveguide Crossing" sch_x=226 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7495 N$29408 N$29410 N$29209 N$29211 "Waveguide Crossing" sch_x=226 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7496 N$29412 N$29414 N$29213 N$29215 "Waveguide Crossing" sch_x=226 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7497 N$29416 N$29418 N$29217 N$29219 "Waveguide Crossing" sch_x=226 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7498 N$29420 N$29422 N$29221 N$29223 "Waveguide Crossing" sch_x=226 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7499 N$29424 N$29426 N$29225 N$29227 "Waveguide Crossing" sch_x=226 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7500 N$29428 N$29430 N$29229 N$29231 "Waveguide Crossing" sch_x=226 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7501 N$29432 N$29434 N$29233 N$29235 "Waveguide Crossing" sch_x=226 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7502 N$29436 N$29438 N$29237 N$29239 "Waveguide Crossing" sch_x=226 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7503 N$29440 N$29442 N$29241 N$29243 "Waveguide Crossing" sch_x=226 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7504 N$29444 N$29446 N$29245 N$29247 "Waveguide Crossing" sch_x=226 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7505 N$29448 N$29450 N$29249 N$29251 "Waveguide Crossing" sch_x=226 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7506 N$29452 N$29454 N$29253 N$29255 "Waveguide Crossing" sch_x=226 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7507 N$29456 N$29458 N$29257 N$29259 "Waveguide Crossing" sch_x=226 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7508 N$29460 N$29462 N$29261 N$29263 "Waveguide Crossing" sch_x=226 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7509 N$29464 N$29466 N$29265 N$29267 "Waveguide Crossing" sch_x=226 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7510 N$29468 N$29470 N$29269 N$29271 "Waveguide Crossing" sch_x=226 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7511 N$29472 N$29474 N$29273 N$29275 "Waveguide Crossing" sch_x=226 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7512 N$29476 N$29478 N$29277 N$29279 "Waveguide Crossing" sch_x=226 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7513 N$29480 N$29482 N$29281 N$29283 "Waveguide Crossing" sch_x=226 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7514 N$29484 N$29486 N$29285 N$29287 "Waveguide Crossing" sch_x=226 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7515 N$29488 N$29490 N$29289 N$29291 "Waveguide Crossing" sch_x=226 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7516 N$29492 N$29494 N$29293 N$29295 "Waveguide Crossing" sch_x=226 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7517 N$29496 N$29498 N$29297 N$29299 "Waveguide Crossing" sch_x=226 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7518 N$29500 N$29502 N$29301 N$29303 "Waveguide Crossing" sch_x=226 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7519 N$29504 N$29506 N$29305 N$29307 "Waveguide Crossing" sch_x=226 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7520 N$29508 N$29510 N$29309 N$29311 "Waveguide Crossing" sch_x=226 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7521 N$29512 N$29514 N$29313 N$29315 "Waveguide Crossing" sch_x=226 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7522 N$29516 N$29518 N$29317 N$29319 "Waveguide Crossing" sch_x=226 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7523 N$29520 N$29522 N$29321 N$29323 "Waveguide Crossing" sch_x=226 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7524 N$29524 N$29526 N$29325 N$29327 "Waveguide Crossing" sch_x=226 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7525 N$29528 N$29530 N$29329 N$29331 "Waveguide Crossing" sch_x=226 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7526 N$29532 N$29534 N$29333 N$29335 "Waveguide Crossing" sch_x=226 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7527 N$29536 N$29538 N$29337 N$29339 "Waveguide Crossing" sch_x=226 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7528 N$29540 N$29542 N$29341 N$29343 "Waveguide Crossing" sch_x=226 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7529 N$29544 N$29546 N$29345 N$29347 "Waveguide Crossing" sch_x=226 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7530 N$29548 N$29550 N$29349 N$29351 "Waveguide Crossing" sch_x=226 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7531 N$29552 N$29554 N$29353 N$29355 "Waveguide Crossing" sch_x=226 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7532 N$29556 N$29558 N$29357 N$29359 "Waveguide Crossing" sch_x=226 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7533 N$29560 N$29562 N$29361 N$29363 "Waveguide Crossing" sch_x=226 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7534 N$29564 N$29566 N$29365 N$29367 "Waveguide Crossing" sch_x=226 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7535 N$29568 N$29570 N$29369 N$29371 "Waveguide Crossing" sch_x=226 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7536 N$29572 N$29574 N$29373 N$29375 "Waveguide Crossing" sch_x=226 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7537 N$29576 N$29578 N$29377 N$29379 "Waveguide Crossing" sch_x=226 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7538 N$29580 N$29582 N$29381 N$29383 "Waveguide Crossing" sch_x=226 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7539 N$29584 N$29586 N$29385 N$29387 "Waveguide Crossing" sch_x=226 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7540 N$29588 N$29590 N$29389 N$29391 "Waveguide Crossing" sch_x=226 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7541 N$29592 N$29594 N$29393 N$29395 "Waveguide Crossing" sch_x=226 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7542 N$29596 N$29598 N$29397 N$29399 "Waveguide Crossing" sch_x=226 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7543 N$29600 N$34529 N$29401 N$29403 "Waveguide Crossing" sch_x=226 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7544 N$34333 N$29602 N$29405 N$29407 "Waveguide Crossing" sch_x=224 sch_y=48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7545 N$29604 N$29606 N$29409 N$29411 "Waveguide Crossing" sch_x=224 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7546 N$29608 N$29610 N$29413 N$29415 "Waveguide Crossing" sch_x=224 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7547 N$29612 N$29614 N$29417 N$29419 "Waveguide Crossing" sch_x=224 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7548 N$29616 N$29618 N$29421 N$29423 "Waveguide Crossing" sch_x=224 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7549 N$29620 N$29622 N$29425 N$29427 "Waveguide Crossing" sch_x=224 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7550 N$29624 N$29626 N$29429 N$29431 "Waveguide Crossing" sch_x=224 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7551 N$29628 N$29630 N$29433 N$29435 "Waveguide Crossing" sch_x=224 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7552 N$29632 N$29634 N$29437 N$29439 "Waveguide Crossing" sch_x=224 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7553 N$29636 N$29638 N$29441 N$29443 "Waveguide Crossing" sch_x=224 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7554 N$29640 N$29642 N$29445 N$29447 "Waveguide Crossing" sch_x=224 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7555 N$29644 N$29646 N$29449 N$29451 "Waveguide Crossing" sch_x=224 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7556 N$29648 N$29650 N$29453 N$29455 "Waveguide Crossing" sch_x=224 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7557 N$29652 N$29654 N$29457 N$29459 "Waveguide Crossing" sch_x=224 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7558 N$29656 N$29658 N$29461 N$29463 "Waveguide Crossing" sch_x=224 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7559 N$29660 N$29662 N$29465 N$29467 "Waveguide Crossing" sch_x=224 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7560 N$29664 N$29666 N$29469 N$29471 "Waveguide Crossing" sch_x=224 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7561 N$29668 N$29670 N$29473 N$29475 "Waveguide Crossing" sch_x=224 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7562 N$29672 N$29674 N$29477 N$29479 "Waveguide Crossing" sch_x=224 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7563 N$29676 N$29678 N$29481 N$29483 "Waveguide Crossing" sch_x=224 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7564 N$29680 N$29682 N$29485 N$29487 "Waveguide Crossing" sch_x=224 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7565 N$29684 N$29686 N$29489 N$29491 "Waveguide Crossing" sch_x=224 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7566 N$29688 N$29690 N$29493 N$29495 "Waveguide Crossing" sch_x=224 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7567 N$29692 N$29694 N$29497 N$29499 "Waveguide Crossing" sch_x=224 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7568 N$29696 N$29698 N$29501 N$29503 "Waveguide Crossing" sch_x=224 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7569 N$29700 N$29702 N$29505 N$29507 "Waveguide Crossing" sch_x=224 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7570 N$29704 N$29706 N$29509 N$29511 "Waveguide Crossing" sch_x=224 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7571 N$29708 N$29710 N$29513 N$29515 "Waveguide Crossing" sch_x=224 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7572 N$29712 N$29714 N$29517 N$29519 "Waveguide Crossing" sch_x=224 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7573 N$29716 N$29718 N$29521 N$29523 "Waveguide Crossing" sch_x=224 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7574 N$29720 N$29722 N$29525 N$29527 "Waveguide Crossing" sch_x=224 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7575 N$29724 N$29726 N$29529 N$29531 "Waveguide Crossing" sch_x=224 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7576 N$29728 N$29730 N$29533 N$29535 "Waveguide Crossing" sch_x=224 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7577 N$29732 N$29734 N$29537 N$29539 "Waveguide Crossing" sch_x=224 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7578 N$29736 N$29738 N$29541 N$29543 "Waveguide Crossing" sch_x=224 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7579 N$29740 N$29742 N$29545 N$29547 "Waveguide Crossing" sch_x=224 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7580 N$29744 N$29746 N$29549 N$29551 "Waveguide Crossing" sch_x=224 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7581 N$29748 N$29750 N$29553 N$29555 "Waveguide Crossing" sch_x=224 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7582 N$29752 N$29754 N$29557 N$29559 "Waveguide Crossing" sch_x=224 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7583 N$29756 N$29758 N$29561 N$29563 "Waveguide Crossing" sch_x=224 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7584 N$29760 N$29762 N$29565 N$29567 "Waveguide Crossing" sch_x=224 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7585 N$29764 N$29766 N$29569 N$29571 "Waveguide Crossing" sch_x=224 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7586 N$29768 N$29770 N$29573 N$29575 "Waveguide Crossing" sch_x=224 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7587 N$29772 N$29774 N$29577 N$29579 "Waveguide Crossing" sch_x=224 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7588 N$29776 N$29778 N$29581 N$29583 "Waveguide Crossing" sch_x=224 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7589 N$29780 N$29782 N$29585 N$29587 "Waveguide Crossing" sch_x=224 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7590 N$29784 N$29786 N$29589 N$29591 "Waveguide Crossing" sch_x=224 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7591 N$29788 N$29790 N$29593 N$29595 "Waveguide Crossing" sch_x=224 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7592 N$29792 N$34527 N$29597 N$29599 "Waveguide Crossing" sch_x=224 sch_y=-48 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7593 N$34335 N$29794 N$29601 N$29603 "Waveguide Crossing" sch_x=222 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7594 N$29796 N$29798 N$29605 N$29607 "Waveguide Crossing" sch_x=222 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7595 N$29800 N$29802 N$29609 N$29611 "Waveguide Crossing" sch_x=222 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7596 N$29804 N$29806 N$29613 N$29615 "Waveguide Crossing" sch_x=222 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7597 N$29808 N$29810 N$29617 N$29619 "Waveguide Crossing" sch_x=222 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7598 N$29812 N$29814 N$29621 N$29623 "Waveguide Crossing" sch_x=222 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7599 N$29816 N$29818 N$29625 N$29627 "Waveguide Crossing" sch_x=222 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7600 N$29820 N$29822 N$29629 N$29631 "Waveguide Crossing" sch_x=222 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7601 N$29824 N$29826 N$29633 N$29635 "Waveguide Crossing" sch_x=222 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7602 N$29828 N$29830 N$29637 N$29639 "Waveguide Crossing" sch_x=222 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7603 N$29832 N$29834 N$29641 N$29643 "Waveguide Crossing" sch_x=222 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7604 N$29836 N$29838 N$29645 N$29647 "Waveguide Crossing" sch_x=222 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7605 N$29840 N$29842 N$29649 N$29651 "Waveguide Crossing" sch_x=222 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7606 N$29844 N$29846 N$29653 N$29655 "Waveguide Crossing" sch_x=222 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7607 N$29848 N$29850 N$29657 N$29659 "Waveguide Crossing" sch_x=222 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7608 N$29852 N$29854 N$29661 N$29663 "Waveguide Crossing" sch_x=222 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7609 N$29856 N$29858 N$29665 N$29667 "Waveguide Crossing" sch_x=222 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7610 N$29860 N$29862 N$29669 N$29671 "Waveguide Crossing" sch_x=222 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7611 N$29864 N$29866 N$29673 N$29675 "Waveguide Crossing" sch_x=222 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7612 N$29868 N$29870 N$29677 N$29679 "Waveguide Crossing" sch_x=222 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7613 N$29872 N$29874 N$29681 N$29683 "Waveguide Crossing" sch_x=222 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7614 N$29876 N$29878 N$29685 N$29687 "Waveguide Crossing" sch_x=222 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7615 N$29880 N$29882 N$29689 N$29691 "Waveguide Crossing" sch_x=222 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7616 N$29884 N$29886 N$29693 N$29695 "Waveguide Crossing" sch_x=222 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7617 N$29888 N$29890 N$29697 N$29699 "Waveguide Crossing" sch_x=222 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7618 N$29892 N$29894 N$29701 N$29703 "Waveguide Crossing" sch_x=222 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7619 N$29896 N$29898 N$29705 N$29707 "Waveguide Crossing" sch_x=222 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7620 N$29900 N$29902 N$29709 N$29711 "Waveguide Crossing" sch_x=222 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7621 N$29904 N$29906 N$29713 N$29715 "Waveguide Crossing" sch_x=222 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7622 N$29908 N$29910 N$29717 N$29719 "Waveguide Crossing" sch_x=222 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7623 N$29912 N$29914 N$29721 N$29723 "Waveguide Crossing" sch_x=222 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7624 N$29916 N$29918 N$29725 N$29727 "Waveguide Crossing" sch_x=222 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7625 N$29920 N$29922 N$29729 N$29731 "Waveguide Crossing" sch_x=222 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7626 N$29924 N$29926 N$29733 N$29735 "Waveguide Crossing" sch_x=222 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7627 N$29928 N$29930 N$29737 N$29739 "Waveguide Crossing" sch_x=222 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7628 N$29932 N$29934 N$29741 N$29743 "Waveguide Crossing" sch_x=222 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7629 N$29936 N$29938 N$29745 N$29747 "Waveguide Crossing" sch_x=222 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7630 N$29940 N$29942 N$29749 N$29751 "Waveguide Crossing" sch_x=222 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7631 N$29944 N$29946 N$29753 N$29755 "Waveguide Crossing" sch_x=222 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7632 N$29948 N$29950 N$29757 N$29759 "Waveguide Crossing" sch_x=222 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7633 N$29952 N$29954 N$29761 N$29763 "Waveguide Crossing" sch_x=222 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7634 N$29956 N$29958 N$29765 N$29767 "Waveguide Crossing" sch_x=222 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7635 N$29960 N$29962 N$29769 N$29771 "Waveguide Crossing" sch_x=222 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7636 N$29964 N$29966 N$29773 N$29775 "Waveguide Crossing" sch_x=222 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7637 N$29968 N$29970 N$29777 N$29779 "Waveguide Crossing" sch_x=222 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7638 N$29972 N$29974 N$29781 N$29783 "Waveguide Crossing" sch_x=222 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7639 N$29976 N$29978 N$29785 N$29787 "Waveguide Crossing" sch_x=222 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7640 N$29980 N$34525 N$29789 N$29791 "Waveguide Crossing" sch_x=222 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7641 N$34337 N$29982 N$29793 N$29795 "Waveguide Crossing" sch_x=220 sch_y=46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7642 N$29984 N$29986 N$29797 N$29799 "Waveguide Crossing" sch_x=220 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7643 N$29988 N$29990 N$29801 N$29803 "Waveguide Crossing" sch_x=220 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7644 N$29992 N$29994 N$29805 N$29807 "Waveguide Crossing" sch_x=220 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7645 N$29996 N$29998 N$29809 N$29811 "Waveguide Crossing" sch_x=220 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7646 N$30000 N$30002 N$29813 N$29815 "Waveguide Crossing" sch_x=220 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7647 N$30004 N$30006 N$29817 N$29819 "Waveguide Crossing" sch_x=220 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7648 N$30008 N$30010 N$29821 N$29823 "Waveguide Crossing" sch_x=220 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7649 N$30012 N$30014 N$29825 N$29827 "Waveguide Crossing" sch_x=220 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7650 N$30016 N$30018 N$29829 N$29831 "Waveguide Crossing" sch_x=220 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7651 N$30020 N$30022 N$29833 N$29835 "Waveguide Crossing" sch_x=220 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7652 N$30024 N$30026 N$29837 N$29839 "Waveguide Crossing" sch_x=220 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7653 N$30028 N$30030 N$29841 N$29843 "Waveguide Crossing" sch_x=220 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7654 N$30032 N$30034 N$29845 N$29847 "Waveguide Crossing" sch_x=220 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7655 N$30036 N$30038 N$29849 N$29851 "Waveguide Crossing" sch_x=220 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7656 N$30040 N$30042 N$29853 N$29855 "Waveguide Crossing" sch_x=220 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7657 N$30044 N$30046 N$29857 N$29859 "Waveguide Crossing" sch_x=220 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7658 N$30048 N$30050 N$29861 N$29863 "Waveguide Crossing" sch_x=220 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7659 N$30052 N$30054 N$29865 N$29867 "Waveguide Crossing" sch_x=220 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7660 N$30056 N$30058 N$29869 N$29871 "Waveguide Crossing" sch_x=220 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7661 N$30060 N$30062 N$29873 N$29875 "Waveguide Crossing" sch_x=220 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7662 N$30064 N$30066 N$29877 N$29879 "Waveguide Crossing" sch_x=220 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7663 N$30068 N$30070 N$29881 N$29883 "Waveguide Crossing" sch_x=220 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7664 N$30072 N$30074 N$29885 N$29887 "Waveguide Crossing" sch_x=220 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7665 N$30076 N$30078 N$29889 N$29891 "Waveguide Crossing" sch_x=220 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7666 N$30080 N$30082 N$29893 N$29895 "Waveguide Crossing" sch_x=220 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7667 N$30084 N$30086 N$29897 N$29899 "Waveguide Crossing" sch_x=220 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7668 N$30088 N$30090 N$29901 N$29903 "Waveguide Crossing" sch_x=220 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7669 N$30092 N$30094 N$29905 N$29907 "Waveguide Crossing" sch_x=220 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7670 N$30096 N$30098 N$29909 N$29911 "Waveguide Crossing" sch_x=220 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7671 N$30100 N$30102 N$29913 N$29915 "Waveguide Crossing" sch_x=220 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7672 N$30104 N$30106 N$29917 N$29919 "Waveguide Crossing" sch_x=220 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7673 N$30108 N$30110 N$29921 N$29923 "Waveguide Crossing" sch_x=220 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7674 N$30112 N$30114 N$29925 N$29927 "Waveguide Crossing" sch_x=220 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7675 N$30116 N$30118 N$29929 N$29931 "Waveguide Crossing" sch_x=220 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7676 N$30120 N$30122 N$29933 N$29935 "Waveguide Crossing" sch_x=220 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7677 N$30124 N$30126 N$29937 N$29939 "Waveguide Crossing" sch_x=220 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7678 N$30128 N$30130 N$29941 N$29943 "Waveguide Crossing" sch_x=220 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7679 N$30132 N$30134 N$29945 N$29947 "Waveguide Crossing" sch_x=220 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7680 N$30136 N$30138 N$29949 N$29951 "Waveguide Crossing" sch_x=220 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7681 N$30140 N$30142 N$29953 N$29955 "Waveguide Crossing" sch_x=220 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7682 N$30144 N$30146 N$29957 N$29959 "Waveguide Crossing" sch_x=220 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7683 N$30148 N$30150 N$29961 N$29963 "Waveguide Crossing" sch_x=220 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7684 N$30152 N$30154 N$29965 N$29967 "Waveguide Crossing" sch_x=220 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7685 N$30156 N$30158 N$29969 N$29971 "Waveguide Crossing" sch_x=220 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7686 N$30160 N$30162 N$29973 N$29975 "Waveguide Crossing" sch_x=220 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7687 N$30164 N$34523 N$29977 N$29979 "Waveguide Crossing" sch_x=220 sch_y=-46 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7688 N$34339 N$30166 N$29981 N$29983 "Waveguide Crossing" sch_x=218 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7689 N$30168 N$30170 N$29985 N$29987 "Waveguide Crossing" sch_x=218 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7690 N$30172 N$30174 N$29989 N$29991 "Waveguide Crossing" sch_x=218 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7691 N$30176 N$30178 N$29993 N$29995 "Waveguide Crossing" sch_x=218 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7692 N$30180 N$30182 N$29997 N$29999 "Waveguide Crossing" sch_x=218 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7693 N$30184 N$30186 N$30001 N$30003 "Waveguide Crossing" sch_x=218 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7694 N$30188 N$30190 N$30005 N$30007 "Waveguide Crossing" sch_x=218 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7695 N$30192 N$30194 N$30009 N$30011 "Waveguide Crossing" sch_x=218 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7696 N$30196 N$30198 N$30013 N$30015 "Waveguide Crossing" sch_x=218 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7697 N$30200 N$30202 N$30017 N$30019 "Waveguide Crossing" sch_x=218 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7698 N$30204 N$30206 N$30021 N$30023 "Waveguide Crossing" sch_x=218 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7699 N$30208 N$30210 N$30025 N$30027 "Waveguide Crossing" sch_x=218 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7700 N$30212 N$30214 N$30029 N$30031 "Waveguide Crossing" sch_x=218 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7701 N$30216 N$30218 N$30033 N$30035 "Waveguide Crossing" sch_x=218 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7702 N$30220 N$30222 N$30037 N$30039 "Waveguide Crossing" sch_x=218 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7703 N$30224 N$30226 N$30041 N$30043 "Waveguide Crossing" sch_x=218 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7704 N$30228 N$30230 N$30045 N$30047 "Waveguide Crossing" sch_x=218 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7705 N$30232 N$30234 N$30049 N$30051 "Waveguide Crossing" sch_x=218 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7706 N$30236 N$30238 N$30053 N$30055 "Waveguide Crossing" sch_x=218 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7707 N$30240 N$30242 N$30057 N$30059 "Waveguide Crossing" sch_x=218 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7708 N$30244 N$30246 N$30061 N$30063 "Waveguide Crossing" sch_x=218 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7709 N$30248 N$30250 N$30065 N$30067 "Waveguide Crossing" sch_x=218 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7710 N$30252 N$30254 N$30069 N$30071 "Waveguide Crossing" sch_x=218 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7711 N$30256 N$30258 N$30073 N$30075 "Waveguide Crossing" sch_x=218 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7712 N$30260 N$30262 N$30077 N$30079 "Waveguide Crossing" sch_x=218 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7713 N$30264 N$30266 N$30081 N$30083 "Waveguide Crossing" sch_x=218 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7714 N$30268 N$30270 N$30085 N$30087 "Waveguide Crossing" sch_x=218 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7715 N$30272 N$30274 N$30089 N$30091 "Waveguide Crossing" sch_x=218 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7716 N$30276 N$30278 N$30093 N$30095 "Waveguide Crossing" sch_x=218 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7717 N$30280 N$30282 N$30097 N$30099 "Waveguide Crossing" sch_x=218 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7718 N$30284 N$30286 N$30101 N$30103 "Waveguide Crossing" sch_x=218 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7719 N$30288 N$30290 N$30105 N$30107 "Waveguide Crossing" sch_x=218 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7720 N$30292 N$30294 N$30109 N$30111 "Waveguide Crossing" sch_x=218 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7721 N$30296 N$30298 N$30113 N$30115 "Waveguide Crossing" sch_x=218 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7722 N$30300 N$30302 N$30117 N$30119 "Waveguide Crossing" sch_x=218 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7723 N$30304 N$30306 N$30121 N$30123 "Waveguide Crossing" sch_x=218 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7724 N$30308 N$30310 N$30125 N$30127 "Waveguide Crossing" sch_x=218 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7725 N$30312 N$30314 N$30129 N$30131 "Waveguide Crossing" sch_x=218 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7726 N$30316 N$30318 N$30133 N$30135 "Waveguide Crossing" sch_x=218 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7727 N$30320 N$30322 N$30137 N$30139 "Waveguide Crossing" sch_x=218 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7728 N$30324 N$30326 N$30141 N$30143 "Waveguide Crossing" sch_x=218 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7729 N$30328 N$30330 N$30145 N$30147 "Waveguide Crossing" sch_x=218 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7730 N$30332 N$30334 N$30149 N$30151 "Waveguide Crossing" sch_x=218 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7731 N$30336 N$30338 N$30153 N$30155 "Waveguide Crossing" sch_x=218 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7732 N$30340 N$30342 N$30157 N$30159 "Waveguide Crossing" sch_x=218 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7733 N$30344 N$34521 N$30161 N$30163 "Waveguide Crossing" sch_x=218 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7734 N$34341 N$30346 N$30165 N$30167 "Waveguide Crossing" sch_x=216 sch_y=44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7735 N$30348 N$30350 N$30169 N$30171 "Waveguide Crossing" sch_x=216 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7736 N$30352 N$30354 N$30173 N$30175 "Waveguide Crossing" sch_x=216 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7737 N$30356 N$30358 N$30177 N$30179 "Waveguide Crossing" sch_x=216 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7738 N$30360 N$30362 N$30181 N$30183 "Waveguide Crossing" sch_x=216 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7739 N$30364 N$30366 N$30185 N$30187 "Waveguide Crossing" sch_x=216 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7740 N$30368 N$30370 N$30189 N$30191 "Waveguide Crossing" sch_x=216 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7741 N$30372 N$30374 N$30193 N$30195 "Waveguide Crossing" sch_x=216 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7742 N$30376 N$30378 N$30197 N$30199 "Waveguide Crossing" sch_x=216 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7743 N$30380 N$30382 N$30201 N$30203 "Waveguide Crossing" sch_x=216 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7744 N$30384 N$30386 N$30205 N$30207 "Waveguide Crossing" sch_x=216 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7745 N$30388 N$30390 N$30209 N$30211 "Waveguide Crossing" sch_x=216 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7746 N$30392 N$30394 N$30213 N$30215 "Waveguide Crossing" sch_x=216 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7747 N$30396 N$30398 N$30217 N$30219 "Waveguide Crossing" sch_x=216 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7748 N$30400 N$30402 N$30221 N$30223 "Waveguide Crossing" sch_x=216 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7749 N$30404 N$30406 N$30225 N$30227 "Waveguide Crossing" sch_x=216 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7750 N$30408 N$30410 N$30229 N$30231 "Waveguide Crossing" sch_x=216 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7751 N$30412 N$30414 N$30233 N$30235 "Waveguide Crossing" sch_x=216 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7752 N$30416 N$30418 N$30237 N$30239 "Waveguide Crossing" sch_x=216 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7753 N$30420 N$30422 N$30241 N$30243 "Waveguide Crossing" sch_x=216 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7754 N$30424 N$30426 N$30245 N$30247 "Waveguide Crossing" sch_x=216 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7755 N$30428 N$30430 N$30249 N$30251 "Waveguide Crossing" sch_x=216 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7756 N$30432 N$30434 N$30253 N$30255 "Waveguide Crossing" sch_x=216 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7757 N$30436 N$30438 N$30257 N$30259 "Waveguide Crossing" sch_x=216 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7758 N$30440 N$30442 N$30261 N$30263 "Waveguide Crossing" sch_x=216 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7759 N$30444 N$30446 N$30265 N$30267 "Waveguide Crossing" sch_x=216 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7760 N$30448 N$30450 N$30269 N$30271 "Waveguide Crossing" sch_x=216 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7761 N$30452 N$30454 N$30273 N$30275 "Waveguide Crossing" sch_x=216 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7762 N$30456 N$30458 N$30277 N$30279 "Waveguide Crossing" sch_x=216 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7763 N$30460 N$30462 N$30281 N$30283 "Waveguide Crossing" sch_x=216 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7764 N$30464 N$30466 N$30285 N$30287 "Waveguide Crossing" sch_x=216 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7765 N$30468 N$30470 N$30289 N$30291 "Waveguide Crossing" sch_x=216 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7766 N$30472 N$30474 N$30293 N$30295 "Waveguide Crossing" sch_x=216 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7767 N$30476 N$30478 N$30297 N$30299 "Waveguide Crossing" sch_x=216 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7768 N$30480 N$30482 N$30301 N$30303 "Waveguide Crossing" sch_x=216 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7769 N$30484 N$30486 N$30305 N$30307 "Waveguide Crossing" sch_x=216 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7770 N$30488 N$30490 N$30309 N$30311 "Waveguide Crossing" sch_x=216 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7771 N$30492 N$30494 N$30313 N$30315 "Waveguide Crossing" sch_x=216 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7772 N$30496 N$30498 N$30317 N$30319 "Waveguide Crossing" sch_x=216 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7773 N$30500 N$30502 N$30321 N$30323 "Waveguide Crossing" sch_x=216 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7774 N$30504 N$30506 N$30325 N$30327 "Waveguide Crossing" sch_x=216 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7775 N$30508 N$30510 N$30329 N$30331 "Waveguide Crossing" sch_x=216 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7776 N$30512 N$30514 N$30333 N$30335 "Waveguide Crossing" sch_x=216 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7777 N$30516 N$30518 N$30337 N$30339 "Waveguide Crossing" sch_x=216 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7778 N$30520 N$34519 N$30341 N$30343 "Waveguide Crossing" sch_x=216 sch_y=-44 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7779 N$34343 N$30522 N$30345 N$30347 "Waveguide Crossing" sch_x=214 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7780 N$30524 N$30526 N$30349 N$30351 "Waveguide Crossing" sch_x=214 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7781 N$30528 N$30530 N$30353 N$30355 "Waveguide Crossing" sch_x=214 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7782 N$30532 N$30534 N$30357 N$30359 "Waveguide Crossing" sch_x=214 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7783 N$30536 N$30538 N$30361 N$30363 "Waveguide Crossing" sch_x=214 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7784 N$30540 N$30542 N$30365 N$30367 "Waveguide Crossing" sch_x=214 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7785 N$30544 N$30546 N$30369 N$30371 "Waveguide Crossing" sch_x=214 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7786 N$30548 N$30550 N$30373 N$30375 "Waveguide Crossing" sch_x=214 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7787 N$30552 N$30554 N$30377 N$30379 "Waveguide Crossing" sch_x=214 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7788 N$30556 N$30558 N$30381 N$30383 "Waveguide Crossing" sch_x=214 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7789 N$30560 N$30562 N$30385 N$30387 "Waveguide Crossing" sch_x=214 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7790 N$30564 N$30566 N$30389 N$30391 "Waveguide Crossing" sch_x=214 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7791 N$30568 N$30570 N$30393 N$30395 "Waveguide Crossing" sch_x=214 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7792 N$30572 N$30574 N$30397 N$30399 "Waveguide Crossing" sch_x=214 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7793 N$30576 N$30578 N$30401 N$30403 "Waveguide Crossing" sch_x=214 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7794 N$30580 N$30582 N$30405 N$30407 "Waveguide Crossing" sch_x=214 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7795 N$30584 N$30586 N$30409 N$30411 "Waveguide Crossing" sch_x=214 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7796 N$30588 N$30590 N$30413 N$30415 "Waveguide Crossing" sch_x=214 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7797 N$30592 N$30594 N$30417 N$30419 "Waveguide Crossing" sch_x=214 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7798 N$30596 N$30598 N$30421 N$30423 "Waveguide Crossing" sch_x=214 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7799 N$30600 N$30602 N$30425 N$30427 "Waveguide Crossing" sch_x=214 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7800 N$30604 N$30606 N$30429 N$30431 "Waveguide Crossing" sch_x=214 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7801 N$30608 N$30610 N$30433 N$30435 "Waveguide Crossing" sch_x=214 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7802 N$30612 N$30614 N$30437 N$30439 "Waveguide Crossing" sch_x=214 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7803 N$30616 N$30618 N$30441 N$30443 "Waveguide Crossing" sch_x=214 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7804 N$30620 N$30622 N$30445 N$30447 "Waveguide Crossing" sch_x=214 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7805 N$30624 N$30626 N$30449 N$30451 "Waveguide Crossing" sch_x=214 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7806 N$30628 N$30630 N$30453 N$30455 "Waveguide Crossing" sch_x=214 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7807 N$30632 N$30634 N$30457 N$30459 "Waveguide Crossing" sch_x=214 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7808 N$30636 N$30638 N$30461 N$30463 "Waveguide Crossing" sch_x=214 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7809 N$30640 N$30642 N$30465 N$30467 "Waveguide Crossing" sch_x=214 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7810 N$30644 N$30646 N$30469 N$30471 "Waveguide Crossing" sch_x=214 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7811 N$30648 N$30650 N$30473 N$30475 "Waveguide Crossing" sch_x=214 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7812 N$30652 N$30654 N$30477 N$30479 "Waveguide Crossing" sch_x=214 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7813 N$30656 N$30658 N$30481 N$30483 "Waveguide Crossing" sch_x=214 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7814 N$30660 N$30662 N$30485 N$30487 "Waveguide Crossing" sch_x=214 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7815 N$30664 N$30666 N$30489 N$30491 "Waveguide Crossing" sch_x=214 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7816 N$30668 N$30670 N$30493 N$30495 "Waveguide Crossing" sch_x=214 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7817 N$30672 N$30674 N$30497 N$30499 "Waveguide Crossing" sch_x=214 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7818 N$30676 N$30678 N$30501 N$30503 "Waveguide Crossing" sch_x=214 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7819 N$30680 N$30682 N$30505 N$30507 "Waveguide Crossing" sch_x=214 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7820 N$30684 N$30686 N$30509 N$30511 "Waveguide Crossing" sch_x=214 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7821 N$30688 N$30690 N$30513 N$30515 "Waveguide Crossing" sch_x=214 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7822 N$30692 N$34517 N$30517 N$30519 "Waveguide Crossing" sch_x=214 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7823 N$34345 N$30694 N$30521 N$30523 "Waveguide Crossing" sch_x=212 sch_y=42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7824 N$30696 N$30698 N$30525 N$30527 "Waveguide Crossing" sch_x=212 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7825 N$30700 N$30702 N$30529 N$30531 "Waveguide Crossing" sch_x=212 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7826 N$30704 N$30706 N$30533 N$30535 "Waveguide Crossing" sch_x=212 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7827 N$30708 N$30710 N$30537 N$30539 "Waveguide Crossing" sch_x=212 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7828 N$30712 N$30714 N$30541 N$30543 "Waveguide Crossing" sch_x=212 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7829 N$30716 N$30718 N$30545 N$30547 "Waveguide Crossing" sch_x=212 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7830 N$30720 N$30722 N$30549 N$30551 "Waveguide Crossing" sch_x=212 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7831 N$30724 N$30726 N$30553 N$30555 "Waveguide Crossing" sch_x=212 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7832 N$30728 N$30730 N$30557 N$30559 "Waveguide Crossing" sch_x=212 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7833 N$30732 N$30734 N$30561 N$30563 "Waveguide Crossing" sch_x=212 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7834 N$30736 N$30738 N$30565 N$30567 "Waveguide Crossing" sch_x=212 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7835 N$30740 N$30742 N$30569 N$30571 "Waveguide Crossing" sch_x=212 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7836 N$30744 N$30746 N$30573 N$30575 "Waveguide Crossing" sch_x=212 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7837 N$30748 N$30750 N$30577 N$30579 "Waveguide Crossing" sch_x=212 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7838 N$30752 N$30754 N$30581 N$30583 "Waveguide Crossing" sch_x=212 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7839 N$30756 N$30758 N$30585 N$30587 "Waveguide Crossing" sch_x=212 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7840 N$30760 N$30762 N$30589 N$30591 "Waveguide Crossing" sch_x=212 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7841 N$30764 N$30766 N$30593 N$30595 "Waveguide Crossing" sch_x=212 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7842 N$30768 N$30770 N$30597 N$30599 "Waveguide Crossing" sch_x=212 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7843 N$30772 N$30774 N$30601 N$30603 "Waveguide Crossing" sch_x=212 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7844 N$30776 N$30778 N$30605 N$30607 "Waveguide Crossing" sch_x=212 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7845 N$30780 N$30782 N$30609 N$30611 "Waveguide Crossing" sch_x=212 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7846 N$30784 N$30786 N$30613 N$30615 "Waveguide Crossing" sch_x=212 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7847 N$30788 N$30790 N$30617 N$30619 "Waveguide Crossing" sch_x=212 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7848 N$30792 N$30794 N$30621 N$30623 "Waveguide Crossing" sch_x=212 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7849 N$30796 N$30798 N$30625 N$30627 "Waveguide Crossing" sch_x=212 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7850 N$30800 N$30802 N$30629 N$30631 "Waveguide Crossing" sch_x=212 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7851 N$30804 N$30806 N$30633 N$30635 "Waveguide Crossing" sch_x=212 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7852 N$30808 N$30810 N$30637 N$30639 "Waveguide Crossing" sch_x=212 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7853 N$30812 N$30814 N$30641 N$30643 "Waveguide Crossing" sch_x=212 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7854 N$30816 N$30818 N$30645 N$30647 "Waveguide Crossing" sch_x=212 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7855 N$30820 N$30822 N$30649 N$30651 "Waveguide Crossing" sch_x=212 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7856 N$30824 N$30826 N$30653 N$30655 "Waveguide Crossing" sch_x=212 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7857 N$30828 N$30830 N$30657 N$30659 "Waveguide Crossing" sch_x=212 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7858 N$30832 N$30834 N$30661 N$30663 "Waveguide Crossing" sch_x=212 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7859 N$30836 N$30838 N$30665 N$30667 "Waveguide Crossing" sch_x=212 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7860 N$30840 N$30842 N$30669 N$30671 "Waveguide Crossing" sch_x=212 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7861 N$30844 N$30846 N$30673 N$30675 "Waveguide Crossing" sch_x=212 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7862 N$30848 N$30850 N$30677 N$30679 "Waveguide Crossing" sch_x=212 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7863 N$30852 N$30854 N$30681 N$30683 "Waveguide Crossing" sch_x=212 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7864 N$30856 N$30858 N$30685 N$30687 "Waveguide Crossing" sch_x=212 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7865 N$30860 N$34515 N$30689 N$30691 "Waveguide Crossing" sch_x=212 sch_y=-42 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7866 N$34347 N$30862 N$30693 N$30695 "Waveguide Crossing" sch_x=210 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7867 N$30864 N$30866 N$30697 N$30699 "Waveguide Crossing" sch_x=210 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7868 N$30868 N$30870 N$30701 N$30703 "Waveguide Crossing" sch_x=210 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7869 N$30872 N$30874 N$30705 N$30707 "Waveguide Crossing" sch_x=210 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7870 N$30876 N$30878 N$30709 N$30711 "Waveguide Crossing" sch_x=210 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7871 N$30880 N$30882 N$30713 N$30715 "Waveguide Crossing" sch_x=210 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7872 N$30884 N$30886 N$30717 N$30719 "Waveguide Crossing" sch_x=210 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7873 N$30888 N$30890 N$30721 N$30723 "Waveguide Crossing" sch_x=210 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7874 N$30892 N$30894 N$30725 N$30727 "Waveguide Crossing" sch_x=210 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7875 N$30896 N$30898 N$30729 N$30731 "Waveguide Crossing" sch_x=210 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7876 N$30900 N$30902 N$30733 N$30735 "Waveguide Crossing" sch_x=210 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7877 N$30904 N$30906 N$30737 N$30739 "Waveguide Crossing" sch_x=210 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7878 N$30908 N$30910 N$30741 N$30743 "Waveguide Crossing" sch_x=210 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7879 N$30912 N$30914 N$30745 N$30747 "Waveguide Crossing" sch_x=210 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7880 N$30916 N$30918 N$30749 N$30751 "Waveguide Crossing" sch_x=210 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7881 N$30920 N$30922 N$30753 N$30755 "Waveguide Crossing" sch_x=210 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7882 N$30924 N$30926 N$30757 N$30759 "Waveguide Crossing" sch_x=210 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7883 N$30928 N$30930 N$30761 N$30763 "Waveguide Crossing" sch_x=210 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7884 N$30932 N$30934 N$30765 N$30767 "Waveguide Crossing" sch_x=210 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7885 N$30936 N$30938 N$30769 N$30771 "Waveguide Crossing" sch_x=210 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7886 N$30940 N$30942 N$30773 N$30775 "Waveguide Crossing" sch_x=210 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7887 N$30944 N$30946 N$30777 N$30779 "Waveguide Crossing" sch_x=210 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7888 N$30948 N$30950 N$30781 N$30783 "Waveguide Crossing" sch_x=210 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7889 N$30952 N$30954 N$30785 N$30787 "Waveguide Crossing" sch_x=210 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7890 N$30956 N$30958 N$30789 N$30791 "Waveguide Crossing" sch_x=210 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7891 N$30960 N$30962 N$30793 N$30795 "Waveguide Crossing" sch_x=210 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7892 N$30964 N$30966 N$30797 N$30799 "Waveguide Crossing" sch_x=210 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7893 N$30968 N$30970 N$30801 N$30803 "Waveguide Crossing" sch_x=210 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7894 N$30972 N$30974 N$30805 N$30807 "Waveguide Crossing" sch_x=210 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7895 N$30976 N$30978 N$30809 N$30811 "Waveguide Crossing" sch_x=210 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7896 N$30980 N$30982 N$30813 N$30815 "Waveguide Crossing" sch_x=210 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7897 N$30984 N$30986 N$30817 N$30819 "Waveguide Crossing" sch_x=210 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7898 N$30988 N$30990 N$30821 N$30823 "Waveguide Crossing" sch_x=210 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7899 N$30992 N$30994 N$30825 N$30827 "Waveguide Crossing" sch_x=210 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7900 N$30996 N$30998 N$30829 N$30831 "Waveguide Crossing" sch_x=210 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7901 N$31000 N$31002 N$30833 N$30835 "Waveguide Crossing" sch_x=210 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7902 N$31004 N$31006 N$30837 N$30839 "Waveguide Crossing" sch_x=210 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7903 N$31008 N$31010 N$30841 N$30843 "Waveguide Crossing" sch_x=210 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7904 N$31012 N$31014 N$30845 N$30847 "Waveguide Crossing" sch_x=210 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7905 N$31016 N$31018 N$30849 N$30851 "Waveguide Crossing" sch_x=210 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7906 N$31020 N$31022 N$30853 N$30855 "Waveguide Crossing" sch_x=210 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7907 N$31024 N$34513 N$30857 N$30859 "Waveguide Crossing" sch_x=210 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7908 N$34349 N$31026 N$30861 N$30863 "Waveguide Crossing" sch_x=208 sch_y=40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7909 N$31028 N$31030 N$30865 N$30867 "Waveguide Crossing" sch_x=208 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7910 N$31032 N$31034 N$30869 N$30871 "Waveguide Crossing" sch_x=208 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7911 N$31036 N$31038 N$30873 N$30875 "Waveguide Crossing" sch_x=208 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7912 N$31040 N$31042 N$30877 N$30879 "Waveguide Crossing" sch_x=208 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7913 N$31044 N$31046 N$30881 N$30883 "Waveguide Crossing" sch_x=208 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7914 N$31048 N$31050 N$30885 N$30887 "Waveguide Crossing" sch_x=208 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7915 N$31052 N$31054 N$30889 N$30891 "Waveguide Crossing" sch_x=208 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7916 N$31056 N$31058 N$30893 N$30895 "Waveguide Crossing" sch_x=208 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7917 N$31060 N$31062 N$30897 N$30899 "Waveguide Crossing" sch_x=208 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7918 N$31064 N$31066 N$30901 N$30903 "Waveguide Crossing" sch_x=208 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7919 N$31068 N$31070 N$30905 N$30907 "Waveguide Crossing" sch_x=208 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7920 N$31072 N$31074 N$30909 N$30911 "Waveguide Crossing" sch_x=208 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7921 N$31076 N$31078 N$30913 N$30915 "Waveguide Crossing" sch_x=208 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7922 N$31080 N$31082 N$30917 N$30919 "Waveguide Crossing" sch_x=208 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7923 N$31084 N$31086 N$30921 N$30923 "Waveguide Crossing" sch_x=208 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7924 N$31088 N$31090 N$30925 N$30927 "Waveguide Crossing" sch_x=208 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7925 N$31092 N$31094 N$30929 N$30931 "Waveguide Crossing" sch_x=208 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7926 N$31096 N$31098 N$30933 N$30935 "Waveguide Crossing" sch_x=208 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7927 N$31100 N$31102 N$30937 N$30939 "Waveguide Crossing" sch_x=208 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7928 N$31104 N$31106 N$30941 N$30943 "Waveguide Crossing" sch_x=208 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7929 N$31108 N$31110 N$30945 N$30947 "Waveguide Crossing" sch_x=208 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7930 N$31112 N$31114 N$30949 N$30951 "Waveguide Crossing" sch_x=208 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7931 N$31116 N$31118 N$30953 N$30955 "Waveguide Crossing" sch_x=208 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7932 N$31120 N$31122 N$30957 N$30959 "Waveguide Crossing" sch_x=208 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7933 N$31124 N$31126 N$30961 N$30963 "Waveguide Crossing" sch_x=208 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7934 N$31128 N$31130 N$30965 N$30967 "Waveguide Crossing" sch_x=208 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7935 N$31132 N$31134 N$30969 N$30971 "Waveguide Crossing" sch_x=208 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7936 N$31136 N$31138 N$30973 N$30975 "Waveguide Crossing" sch_x=208 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7937 N$31140 N$31142 N$30977 N$30979 "Waveguide Crossing" sch_x=208 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7938 N$31144 N$31146 N$30981 N$30983 "Waveguide Crossing" sch_x=208 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7939 N$31148 N$31150 N$30985 N$30987 "Waveguide Crossing" sch_x=208 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7940 N$31152 N$31154 N$30989 N$30991 "Waveguide Crossing" sch_x=208 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7941 N$31156 N$31158 N$30993 N$30995 "Waveguide Crossing" sch_x=208 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7942 N$31160 N$31162 N$30997 N$30999 "Waveguide Crossing" sch_x=208 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7943 N$31164 N$31166 N$31001 N$31003 "Waveguide Crossing" sch_x=208 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7944 N$31168 N$31170 N$31005 N$31007 "Waveguide Crossing" sch_x=208 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7945 N$31172 N$31174 N$31009 N$31011 "Waveguide Crossing" sch_x=208 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7946 N$31176 N$31178 N$31013 N$31015 "Waveguide Crossing" sch_x=208 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7947 N$31180 N$31182 N$31017 N$31019 "Waveguide Crossing" sch_x=208 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7948 N$31184 N$34511 N$31021 N$31023 "Waveguide Crossing" sch_x=208 sch_y=-40 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7949 N$34351 N$31186 N$31025 N$31027 "Waveguide Crossing" sch_x=206 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7950 N$31188 N$31190 N$31029 N$31031 "Waveguide Crossing" sch_x=206 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7951 N$31192 N$31194 N$31033 N$31035 "Waveguide Crossing" sch_x=206 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7952 N$31196 N$31198 N$31037 N$31039 "Waveguide Crossing" sch_x=206 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7953 N$31200 N$31202 N$31041 N$31043 "Waveguide Crossing" sch_x=206 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7954 N$31204 N$31206 N$31045 N$31047 "Waveguide Crossing" sch_x=206 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7955 N$31208 N$31210 N$31049 N$31051 "Waveguide Crossing" sch_x=206 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7956 N$31212 N$31214 N$31053 N$31055 "Waveguide Crossing" sch_x=206 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7957 N$31216 N$31218 N$31057 N$31059 "Waveguide Crossing" sch_x=206 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7958 N$31220 N$31222 N$31061 N$31063 "Waveguide Crossing" sch_x=206 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7959 N$31224 N$31226 N$31065 N$31067 "Waveguide Crossing" sch_x=206 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7960 N$31228 N$31230 N$31069 N$31071 "Waveguide Crossing" sch_x=206 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7961 N$31232 N$31234 N$31073 N$31075 "Waveguide Crossing" sch_x=206 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7962 N$31236 N$31238 N$31077 N$31079 "Waveguide Crossing" sch_x=206 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7963 N$31240 N$31242 N$31081 N$31083 "Waveguide Crossing" sch_x=206 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7964 N$31244 N$31246 N$31085 N$31087 "Waveguide Crossing" sch_x=206 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7965 N$31248 N$31250 N$31089 N$31091 "Waveguide Crossing" sch_x=206 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7966 N$31252 N$31254 N$31093 N$31095 "Waveguide Crossing" sch_x=206 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7967 N$31256 N$31258 N$31097 N$31099 "Waveguide Crossing" sch_x=206 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7968 N$31260 N$31262 N$31101 N$31103 "Waveguide Crossing" sch_x=206 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7969 N$31264 N$31266 N$31105 N$31107 "Waveguide Crossing" sch_x=206 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7970 N$31268 N$31270 N$31109 N$31111 "Waveguide Crossing" sch_x=206 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7971 N$31272 N$31274 N$31113 N$31115 "Waveguide Crossing" sch_x=206 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7972 N$31276 N$31278 N$31117 N$31119 "Waveguide Crossing" sch_x=206 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7973 N$31280 N$31282 N$31121 N$31123 "Waveguide Crossing" sch_x=206 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7974 N$31284 N$31286 N$31125 N$31127 "Waveguide Crossing" sch_x=206 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7975 N$31288 N$31290 N$31129 N$31131 "Waveguide Crossing" sch_x=206 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7976 N$31292 N$31294 N$31133 N$31135 "Waveguide Crossing" sch_x=206 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7977 N$31296 N$31298 N$31137 N$31139 "Waveguide Crossing" sch_x=206 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7978 N$31300 N$31302 N$31141 N$31143 "Waveguide Crossing" sch_x=206 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7979 N$31304 N$31306 N$31145 N$31147 "Waveguide Crossing" sch_x=206 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7980 N$31308 N$31310 N$31149 N$31151 "Waveguide Crossing" sch_x=206 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7981 N$31312 N$31314 N$31153 N$31155 "Waveguide Crossing" sch_x=206 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7982 N$31316 N$31318 N$31157 N$31159 "Waveguide Crossing" sch_x=206 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7983 N$31320 N$31322 N$31161 N$31163 "Waveguide Crossing" sch_x=206 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7984 N$31324 N$31326 N$31165 N$31167 "Waveguide Crossing" sch_x=206 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7985 N$31328 N$31330 N$31169 N$31171 "Waveguide Crossing" sch_x=206 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7986 N$31332 N$31334 N$31173 N$31175 "Waveguide Crossing" sch_x=206 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7987 N$31336 N$31338 N$31177 N$31179 "Waveguide Crossing" sch_x=206 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7988 N$31340 N$34509 N$31181 N$31183 "Waveguide Crossing" sch_x=206 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7989 N$34353 N$31342 N$31185 N$31187 "Waveguide Crossing" sch_x=204 sch_y=38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7990 N$31344 N$31346 N$31189 N$31191 "Waveguide Crossing" sch_x=204 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7991 N$31348 N$31350 N$31193 N$31195 "Waveguide Crossing" sch_x=204 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7992 N$31352 N$31354 N$31197 N$31199 "Waveguide Crossing" sch_x=204 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7993 N$31356 N$31358 N$31201 N$31203 "Waveguide Crossing" sch_x=204 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7994 N$31360 N$31362 N$31205 N$31207 "Waveguide Crossing" sch_x=204 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7995 N$31364 N$31366 N$31209 N$31211 "Waveguide Crossing" sch_x=204 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7996 N$31368 N$31370 N$31213 N$31215 "Waveguide Crossing" sch_x=204 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7997 N$31372 N$31374 N$31217 N$31219 "Waveguide Crossing" sch_x=204 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7998 N$31376 N$31378 N$31221 N$31223 "Waveguide Crossing" sch_x=204 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C7999 N$31380 N$31382 N$31225 N$31227 "Waveguide Crossing" sch_x=204 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8000 N$31384 N$31386 N$31229 N$31231 "Waveguide Crossing" sch_x=204 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8001 N$31388 N$31390 N$31233 N$31235 "Waveguide Crossing" sch_x=204 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8002 N$31392 N$31394 N$31237 N$31239 "Waveguide Crossing" sch_x=204 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8003 N$31396 N$31398 N$31241 N$31243 "Waveguide Crossing" sch_x=204 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8004 N$31400 N$31402 N$31245 N$31247 "Waveguide Crossing" sch_x=204 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8005 N$31404 N$31406 N$31249 N$31251 "Waveguide Crossing" sch_x=204 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8006 N$31408 N$31410 N$31253 N$31255 "Waveguide Crossing" sch_x=204 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8007 N$31412 N$31414 N$31257 N$31259 "Waveguide Crossing" sch_x=204 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8008 N$31416 N$31418 N$31261 N$31263 "Waveguide Crossing" sch_x=204 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8009 N$31420 N$31422 N$31265 N$31267 "Waveguide Crossing" sch_x=204 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8010 N$31424 N$31426 N$31269 N$31271 "Waveguide Crossing" sch_x=204 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8011 N$31428 N$31430 N$31273 N$31275 "Waveguide Crossing" sch_x=204 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8012 N$31432 N$31434 N$31277 N$31279 "Waveguide Crossing" sch_x=204 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8013 N$31436 N$31438 N$31281 N$31283 "Waveguide Crossing" sch_x=204 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8014 N$31440 N$31442 N$31285 N$31287 "Waveguide Crossing" sch_x=204 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8015 N$31444 N$31446 N$31289 N$31291 "Waveguide Crossing" sch_x=204 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8016 N$31448 N$31450 N$31293 N$31295 "Waveguide Crossing" sch_x=204 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8017 N$31452 N$31454 N$31297 N$31299 "Waveguide Crossing" sch_x=204 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8018 N$31456 N$31458 N$31301 N$31303 "Waveguide Crossing" sch_x=204 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8019 N$31460 N$31462 N$31305 N$31307 "Waveguide Crossing" sch_x=204 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8020 N$31464 N$31466 N$31309 N$31311 "Waveguide Crossing" sch_x=204 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8021 N$31468 N$31470 N$31313 N$31315 "Waveguide Crossing" sch_x=204 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8022 N$31472 N$31474 N$31317 N$31319 "Waveguide Crossing" sch_x=204 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8023 N$31476 N$31478 N$31321 N$31323 "Waveguide Crossing" sch_x=204 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8024 N$31480 N$31482 N$31325 N$31327 "Waveguide Crossing" sch_x=204 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8025 N$31484 N$31486 N$31329 N$31331 "Waveguide Crossing" sch_x=204 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8026 N$31488 N$31490 N$31333 N$31335 "Waveguide Crossing" sch_x=204 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8027 N$31492 N$34507 N$31337 N$31339 "Waveguide Crossing" sch_x=204 sch_y=-38 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8028 N$34355 N$31494 N$31341 N$31343 "Waveguide Crossing" sch_x=202 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8029 N$31496 N$31498 N$31345 N$31347 "Waveguide Crossing" sch_x=202 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8030 N$31500 N$31502 N$31349 N$31351 "Waveguide Crossing" sch_x=202 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8031 N$31504 N$31506 N$31353 N$31355 "Waveguide Crossing" sch_x=202 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8032 N$31508 N$31510 N$31357 N$31359 "Waveguide Crossing" sch_x=202 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8033 N$31512 N$31514 N$31361 N$31363 "Waveguide Crossing" sch_x=202 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8034 N$31516 N$31518 N$31365 N$31367 "Waveguide Crossing" sch_x=202 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8035 N$31520 N$31522 N$31369 N$31371 "Waveguide Crossing" sch_x=202 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8036 N$31524 N$31526 N$31373 N$31375 "Waveguide Crossing" sch_x=202 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8037 N$31528 N$31530 N$31377 N$31379 "Waveguide Crossing" sch_x=202 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8038 N$31532 N$31534 N$31381 N$31383 "Waveguide Crossing" sch_x=202 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8039 N$31536 N$31538 N$31385 N$31387 "Waveguide Crossing" sch_x=202 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8040 N$31540 N$31542 N$31389 N$31391 "Waveguide Crossing" sch_x=202 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8041 N$31544 N$31546 N$31393 N$31395 "Waveguide Crossing" sch_x=202 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8042 N$31548 N$31550 N$31397 N$31399 "Waveguide Crossing" sch_x=202 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8043 N$31552 N$31554 N$31401 N$31403 "Waveguide Crossing" sch_x=202 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8044 N$31556 N$31558 N$31405 N$31407 "Waveguide Crossing" sch_x=202 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8045 N$31560 N$31562 N$31409 N$31411 "Waveguide Crossing" sch_x=202 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8046 N$31564 N$31566 N$31413 N$31415 "Waveguide Crossing" sch_x=202 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8047 N$31568 N$31570 N$31417 N$31419 "Waveguide Crossing" sch_x=202 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8048 N$31572 N$31574 N$31421 N$31423 "Waveguide Crossing" sch_x=202 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8049 N$31576 N$31578 N$31425 N$31427 "Waveguide Crossing" sch_x=202 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8050 N$31580 N$31582 N$31429 N$31431 "Waveguide Crossing" sch_x=202 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8051 N$31584 N$31586 N$31433 N$31435 "Waveguide Crossing" sch_x=202 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8052 N$31588 N$31590 N$31437 N$31439 "Waveguide Crossing" sch_x=202 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8053 N$31592 N$31594 N$31441 N$31443 "Waveguide Crossing" sch_x=202 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8054 N$31596 N$31598 N$31445 N$31447 "Waveguide Crossing" sch_x=202 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8055 N$31600 N$31602 N$31449 N$31451 "Waveguide Crossing" sch_x=202 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8056 N$31604 N$31606 N$31453 N$31455 "Waveguide Crossing" sch_x=202 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8057 N$31608 N$31610 N$31457 N$31459 "Waveguide Crossing" sch_x=202 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8058 N$31612 N$31614 N$31461 N$31463 "Waveguide Crossing" sch_x=202 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8059 N$31616 N$31618 N$31465 N$31467 "Waveguide Crossing" sch_x=202 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8060 N$31620 N$31622 N$31469 N$31471 "Waveguide Crossing" sch_x=202 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8061 N$31624 N$31626 N$31473 N$31475 "Waveguide Crossing" sch_x=202 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8062 N$31628 N$31630 N$31477 N$31479 "Waveguide Crossing" sch_x=202 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8063 N$31632 N$31634 N$31481 N$31483 "Waveguide Crossing" sch_x=202 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8064 N$31636 N$31638 N$31485 N$31487 "Waveguide Crossing" sch_x=202 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8065 N$31640 N$34505 N$31489 N$31491 "Waveguide Crossing" sch_x=202 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8066 N$34357 N$31642 N$31493 N$31495 "Waveguide Crossing" sch_x=200 sch_y=36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8067 N$31644 N$31646 N$31497 N$31499 "Waveguide Crossing" sch_x=200 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8068 N$31648 N$31650 N$31501 N$31503 "Waveguide Crossing" sch_x=200 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8069 N$31652 N$31654 N$31505 N$31507 "Waveguide Crossing" sch_x=200 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8070 N$31656 N$31658 N$31509 N$31511 "Waveguide Crossing" sch_x=200 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8071 N$31660 N$31662 N$31513 N$31515 "Waveguide Crossing" sch_x=200 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8072 N$31664 N$31666 N$31517 N$31519 "Waveguide Crossing" sch_x=200 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8073 N$31668 N$31670 N$31521 N$31523 "Waveguide Crossing" sch_x=200 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8074 N$31672 N$31674 N$31525 N$31527 "Waveguide Crossing" sch_x=200 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8075 N$31676 N$31678 N$31529 N$31531 "Waveguide Crossing" sch_x=200 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8076 N$31680 N$31682 N$31533 N$31535 "Waveguide Crossing" sch_x=200 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8077 N$31684 N$31686 N$31537 N$31539 "Waveguide Crossing" sch_x=200 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8078 N$31688 N$31690 N$31541 N$31543 "Waveguide Crossing" sch_x=200 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8079 N$31692 N$31694 N$31545 N$31547 "Waveguide Crossing" sch_x=200 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8080 N$31696 N$31698 N$31549 N$31551 "Waveguide Crossing" sch_x=200 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8081 N$31700 N$31702 N$31553 N$31555 "Waveguide Crossing" sch_x=200 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8082 N$31704 N$31706 N$31557 N$31559 "Waveguide Crossing" sch_x=200 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8083 N$31708 N$31710 N$31561 N$31563 "Waveguide Crossing" sch_x=200 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8084 N$31712 N$31714 N$31565 N$31567 "Waveguide Crossing" sch_x=200 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8085 N$31716 N$31718 N$31569 N$31571 "Waveguide Crossing" sch_x=200 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8086 N$31720 N$31722 N$31573 N$31575 "Waveguide Crossing" sch_x=200 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8087 N$31724 N$31726 N$31577 N$31579 "Waveguide Crossing" sch_x=200 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8088 N$31728 N$31730 N$31581 N$31583 "Waveguide Crossing" sch_x=200 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8089 N$31732 N$31734 N$31585 N$31587 "Waveguide Crossing" sch_x=200 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8090 N$31736 N$31738 N$31589 N$31591 "Waveguide Crossing" sch_x=200 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8091 N$31740 N$31742 N$31593 N$31595 "Waveguide Crossing" sch_x=200 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8092 N$31744 N$31746 N$31597 N$31599 "Waveguide Crossing" sch_x=200 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8093 N$31748 N$31750 N$31601 N$31603 "Waveguide Crossing" sch_x=200 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8094 N$31752 N$31754 N$31605 N$31607 "Waveguide Crossing" sch_x=200 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8095 N$31756 N$31758 N$31609 N$31611 "Waveguide Crossing" sch_x=200 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8096 N$31760 N$31762 N$31613 N$31615 "Waveguide Crossing" sch_x=200 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8097 N$31764 N$31766 N$31617 N$31619 "Waveguide Crossing" sch_x=200 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8098 N$31768 N$31770 N$31621 N$31623 "Waveguide Crossing" sch_x=200 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8099 N$31772 N$31774 N$31625 N$31627 "Waveguide Crossing" sch_x=200 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8100 N$31776 N$31778 N$31629 N$31631 "Waveguide Crossing" sch_x=200 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8101 N$31780 N$31782 N$31633 N$31635 "Waveguide Crossing" sch_x=200 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8102 N$31784 N$34503 N$31637 N$31639 "Waveguide Crossing" sch_x=200 sch_y=-36 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8103 N$34359 N$31786 N$31641 N$31643 "Waveguide Crossing" sch_x=198 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8104 N$31788 N$31790 N$31645 N$31647 "Waveguide Crossing" sch_x=198 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8105 N$31792 N$31794 N$31649 N$31651 "Waveguide Crossing" sch_x=198 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8106 N$31796 N$31798 N$31653 N$31655 "Waveguide Crossing" sch_x=198 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8107 N$31800 N$31802 N$31657 N$31659 "Waveguide Crossing" sch_x=198 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8108 N$31804 N$31806 N$31661 N$31663 "Waveguide Crossing" sch_x=198 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8109 N$31808 N$31810 N$31665 N$31667 "Waveguide Crossing" sch_x=198 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8110 N$31812 N$31814 N$31669 N$31671 "Waveguide Crossing" sch_x=198 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8111 N$31816 N$31818 N$31673 N$31675 "Waveguide Crossing" sch_x=198 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8112 N$31820 N$31822 N$31677 N$31679 "Waveguide Crossing" sch_x=198 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8113 N$31824 N$31826 N$31681 N$31683 "Waveguide Crossing" sch_x=198 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8114 N$31828 N$31830 N$31685 N$31687 "Waveguide Crossing" sch_x=198 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8115 N$31832 N$31834 N$31689 N$31691 "Waveguide Crossing" sch_x=198 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8116 N$31836 N$31838 N$31693 N$31695 "Waveguide Crossing" sch_x=198 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8117 N$31840 N$31842 N$31697 N$31699 "Waveguide Crossing" sch_x=198 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8118 N$31844 N$31846 N$31701 N$31703 "Waveguide Crossing" sch_x=198 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8119 N$31848 N$31850 N$31705 N$31707 "Waveguide Crossing" sch_x=198 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8120 N$31852 N$31854 N$31709 N$31711 "Waveguide Crossing" sch_x=198 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8121 N$31856 N$31858 N$31713 N$31715 "Waveguide Crossing" sch_x=198 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8122 N$31860 N$31862 N$31717 N$31719 "Waveguide Crossing" sch_x=198 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8123 N$31864 N$31866 N$31721 N$31723 "Waveguide Crossing" sch_x=198 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8124 N$31868 N$31870 N$31725 N$31727 "Waveguide Crossing" sch_x=198 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8125 N$31872 N$31874 N$31729 N$31731 "Waveguide Crossing" sch_x=198 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8126 N$31876 N$31878 N$31733 N$31735 "Waveguide Crossing" sch_x=198 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8127 N$31880 N$31882 N$31737 N$31739 "Waveguide Crossing" sch_x=198 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8128 N$31884 N$31886 N$31741 N$31743 "Waveguide Crossing" sch_x=198 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8129 N$31888 N$31890 N$31745 N$31747 "Waveguide Crossing" sch_x=198 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8130 N$31892 N$31894 N$31749 N$31751 "Waveguide Crossing" sch_x=198 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8131 N$31896 N$31898 N$31753 N$31755 "Waveguide Crossing" sch_x=198 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8132 N$31900 N$31902 N$31757 N$31759 "Waveguide Crossing" sch_x=198 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8133 N$31904 N$31906 N$31761 N$31763 "Waveguide Crossing" sch_x=198 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8134 N$31908 N$31910 N$31765 N$31767 "Waveguide Crossing" sch_x=198 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8135 N$31912 N$31914 N$31769 N$31771 "Waveguide Crossing" sch_x=198 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8136 N$31916 N$31918 N$31773 N$31775 "Waveguide Crossing" sch_x=198 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8137 N$31920 N$31922 N$31777 N$31779 "Waveguide Crossing" sch_x=198 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8138 N$31924 N$34501 N$31781 N$31783 "Waveguide Crossing" sch_x=198 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8139 N$34361 N$31926 N$31785 N$31787 "Waveguide Crossing" sch_x=196 sch_y=34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8140 N$31928 N$31930 N$31789 N$31791 "Waveguide Crossing" sch_x=196 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8141 N$31932 N$31934 N$31793 N$31795 "Waveguide Crossing" sch_x=196 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8142 N$31936 N$31938 N$31797 N$31799 "Waveguide Crossing" sch_x=196 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8143 N$31940 N$31942 N$31801 N$31803 "Waveguide Crossing" sch_x=196 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8144 N$31944 N$31946 N$31805 N$31807 "Waveguide Crossing" sch_x=196 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8145 N$31948 N$31950 N$31809 N$31811 "Waveguide Crossing" sch_x=196 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8146 N$31952 N$31954 N$31813 N$31815 "Waveguide Crossing" sch_x=196 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8147 N$31956 N$31958 N$31817 N$31819 "Waveguide Crossing" sch_x=196 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8148 N$31960 N$31962 N$31821 N$31823 "Waveguide Crossing" sch_x=196 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8149 N$31964 N$31966 N$31825 N$31827 "Waveguide Crossing" sch_x=196 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8150 N$31968 N$31970 N$31829 N$31831 "Waveguide Crossing" sch_x=196 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8151 N$31972 N$31974 N$31833 N$31835 "Waveguide Crossing" sch_x=196 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8152 N$31976 N$31978 N$31837 N$31839 "Waveguide Crossing" sch_x=196 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8153 N$31980 N$31982 N$31841 N$31843 "Waveguide Crossing" sch_x=196 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8154 N$31984 N$31986 N$31845 N$31847 "Waveguide Crossing" sch_x=196 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8155 N$31988 N$31990 N$31849 N$31851 "Waveguide Crossing" sch_x=196 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8156 N$31992 N$31994 N$31853 N$31855 "Waveguide Crossing" sch_x=196 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8157 N$31996 N$31998 N$31857 N$31859 "Waveguide Crossing" sch_x=196 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8158 N$32000 N$32002 N$31861 N$31863 "Waveguide Crossing" sch_x=196 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8159 N$32004 N$32006 N$31865 N$31867 "Waveguide Crossing" sch_x=196 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8160 N$32008 N$32010 N$31869 N$31871 "Waveguide Crossing" sch_x=196 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8161 N$32012 N$32014 N$31873 N$31875 "Waveguide Crossing" sch_x=196 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8162 N$32016 N$32018 N$31877 N$31879 "Waveguide Crossing" sch_x=196 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8163 N$32020 N$32022 N$31881 N$31883 "Waveguide Crossing" sch_x=196 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8164 N$32024 N$32026 N$31885 N$31887 "Waveguide Crossing" sch_x=196 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8165 N$32028 N$32030 N$31889 N$31891 "Waveguide Crossing" sch_x=196 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8166 N$32032 N$32034 N$31893 N$31895 "Waveguide Crossing" sch_x=196 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8167 N$32036 N$32038 N$31897 N$31899 "Waveguide Crossing" sch_x=196 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8168 N$32040 N$32042 N$31901 N$31903 "Waveguide Crossing" sch_x=196 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8169 N$32044 N$32046 N$31905 N$31907 "Waveguide Crossing" sch_x=196 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8170 N$32048 N$32050 N$31909 N$31911 "Waveguide Crossing" sch_x=196 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8171 N$32052 N$32054 N$31913 N$31915 "Waveguide Crossing" sch_x=196 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8172 N$32056 N$32058 N$31917 N$31919 "Waveguide Crossing" sch_x=196 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8173 N$32060 N$34499 N$31921 N$31923 "Waveguide Crossing" sch_x=196 sch_y=-34 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8174 N$34363 N$32062 N$31925 N$31927 "Waveguide Crossing" sch_x=194 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8175 N$32064 N$32066 N$31929 N$31931 "Waveguide Crossing" sch_x=194 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8176 N$32068 N$32070 N$31933 N$31935 "Waveguide Crossing" sch_x=194 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8177 N$32072 N$32074 N$31937 N$31939 "Waveguide Crossing" sch_x=194 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8178 N$32076 N$32078 N$31941 N$31943 "Waveguide Crossing" sch_x=194 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8179 N$32080 N$32082 N$31945 N$31947 "Waveguide Crossing" sch_x=194 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8180 N$32084 N$32086 N$31949 N$31951 "Waveguide Crossing" sch_x=194 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8181 N$32088 N$32090 N$31953 N$31955 "Waveguide Crossing" sch_x=194 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8182 N$32092 N$32094 N$31957 N$31959 "Waveguide Crossing" sch_x=194 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8183 N$32096 N$32098 N$31961 N$31963 "Waveguide Crossing" sch_x=194 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8184 N$32100 N$32102 N$31965 N$31967 "Waveguide Crossing" sch_x=194 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8185 N$32104 N$32106 N$31969 N$31971 "Waveguide Crossing" sch_x=194 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8186 N$32108 N$32110 N$31973 N$31975 "Waveguide Crossing" sch_x=194 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8187 N$32112 N$32114 N$31977 N$31979 "Waveguide Crossing" sch_x=194 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8188 N$32116 N$32118 N$31981 N$31983 "Waveguide Crossing" sch_x=194 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8189 N$32120 N$32122 N$31985 N$31987 "Waveguide Crossing" sch_x=194 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8190 N$32124 N$32126 N$31989 N$31991 "Waveguide Crossing" sch_x=194 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8191 N$32128 N$32130 N$31993 N$31995 "Waveguide Crossing" sch_x=194 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8192 N$32132 N$32134 N$31997 N$31999 "Waveguide Crossing" sch_x=194 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8193 N$32136 N$32138 N$32001 N$32003 "Waveguide Crossing" sch_x=194 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8194 N$32140 N$32142 N$32005 N$32007 "Waveguide Crossing" sch_x=194 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8195 N$32144 N$32146 N$32009 N$32011 "Waveguide Crossing" sch_x=194 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8196 N$32148 N$32150 N$32013 N$32015 "Waveguide Crossing" sch_x=194 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8197 N$32152 N$32154 N$32017 N$32019 "Waveguide Crossing" sch_x=194 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8198 N$32156 N$32158 N$32021 N$32023 "Waveguide Crossing" sch_x=194 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8199 N$32160 N$32162 N$32025 N$32027 "Waveguide Crossing" sch_x=194 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8200 N$32164 N$32166 N$32029 N$32031 "Waveguide Crossing" sch_x=194 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8201 N$32168 N$32170 N$32033 N$32035 "Waveguide Crossing" sch_x=194 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8202 N$32172 N$32174 N$32037 N$32039 "Waveguide Crossing" sch_x=194 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8203 N$32176 N$32178 N$32041 N$32043 "Waveguide Crossing" sch_x=194 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8204 N$32180 N$32182 N$32045 N$32047 "Waveguide Crossing" sch_x=194 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8205 N$32184 N$32186 N$32049 N$32051 "Waveguide Crossing" sch_x=194 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8206 N$32188 N$32190 N$32053 N$32055 "Waveguide Crossing" sch_x=194 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8207 N$32192 N$34497 N$32057 N$32059 "Waveguide Crossing" sch_x=194 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8208 N$34365 N$32194 N$32061 N$32063 "Waveguide Crossing" sch_x=192 sch_y=32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8209 N$32196 N$32198 N$32065 N$32067 "Waveguide Crossing" sch_x=192 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8210 N$32200 N$32202 N$32069 N$32071 "Waveguide Crossing" sch_x=192 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8211 N$32204 N$32206 N$32073 N$32075 "Waveguide Crossing" sch_x=192 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8212 N$32208 N$32210 N$32077 N$32079 "Waveguide Crossing" sch_x=192 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8213 N$32212 N$32214 N$32081 N$32083 "Waveguide Crossing" sch_x=192 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8214 N$32216 N$32218 N$32085 N$32087 "Waveguide Crossing" sch_x=192 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8215 N$32220 N$32222 N$32089 N$32091 "Waveguide Crossing" sch_x=192 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8216 N$32224 N$32226 N$32093 N$32095 "Waveguide Crossing" sch_x=192 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8217 N$32228 N$32230 N$32097 N$32099 "Waveguide Crossing" sch_x=192 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8218 N$32232 N$32234 N$32101 N$32103 "Waveguide Crossing" sch_x=192 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8219 N$32236 N$32238 N$32105 N$32107 "Waveguide Crossing" sch_x=192 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8220 N$32240 N$32242 N$32109 N$32111 "Waveguide Crossing" sch_x=192 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8221 N$32244 N$32246 N$32113 N$32115 "Waveguide Crossing" sch_x=192 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8222 N$32248 N$32250 N$32117 N$32119 "Waveguide Crossing" sch_x=192 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8223 N$32252 N$32254 N$32121 N$32123 "Waveguide Crossing" sch_x=192 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8224 N$32256 N$32258 N$32125 N$32127 "Waveguide Crossing" sch_x=192 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8225 N$32260 N$32262 N$32129 N$32131 "Waveguide Crossing" sch_x=192 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8226 N$32264 N$32266 N$32133 N$32135 "Waveguide Crossing" sch_x=192 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8227 N$32268 N$32270 N$32137 N$32139 "Waveguide Crossing" sch_x=192 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8228 N$32272 N$32274 N$32141 N$32143 "Waveguide Crossing" sch_x=192 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8229 N$32276 N$32278 N$32145 N$32147 "Waveguide Crossing" sch_x=192 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8230 N$32280 N$32282 N$32149 N$32151 "Waveguide Crossing" sch_x=192 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8231 N$32284 N$32286 N$32153 N$32155 "Waveguide Crossing" sch_x=192 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8232 N$32288 N$32290 N$32157 N$32159 "Waveguide Crossing" sch_x=192 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8233 N$32292 N$32294 N$32161 N$32163 "Waveguide Crossing" sch_x=192 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8234 N$32296 N$32298 N$32165 N$32167 "Waveguide Crossing" sch_x=192 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8235 N$32300 N$32302 N$32169 N$32171 "Waveguide Crossing" sch_x=192 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8236 N$32304 N$32306 N$32173 N$32175 "Waveguide Crossing" sch_x=192 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8237 N$32308 N$32310 N$32177 N$32179 "Waveguide Crossing" sch_x=192 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8238 N$32312 N$32314 N$32181 N$32183 "Waveguide Crossing" sch_x=192 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8239 N$32316 N$32318 N$32185 N$32187 "Waveguide Crossing" sch_x=192 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8240 N$32320 N$34495 N$32189 N$32191 "Waveguide Crossing" sch_x=192 sch_y=-32 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8241 N$34367 N$32322 N$32193 N$32195 "Waveguide Crossing" sch_x=190 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8242 N$32324 N$32326 N$32197 N$32199 "Waveguide Crossing" sch_x=190 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8243 N$32328 N$32330 N$32201 N$32203 "Waveguide Crossing" sch_x=190 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8244 N$32332 N$32334 N$32205 N$32207 "Waveguide Crossing" sch_x=190 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8245 N$32336 N$32338 N$32209 N$32211 "Waveguide Crossing" sch_x=190 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8246 N$32340 N$32342 N$32213 N$32215 "Waveguide Crossing" sch_x=190 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8247 N$32344 N$32346 N$32217 N$32219 "Waveguide Crossing" sch_x=190 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8248 N$32348 N$32350 N$32221 N$32223 "Waveguide Crossing" sch_x=190 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8249 N$32352 N$32354 N$32225 N$32227 "Waveguide Crossing" sch_x=190 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8250 N$32356 N$32358 N$32229 N$32231 "Waveguide Crossing" sch_x=190 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8251 N$32360 N$32362 N$32233 N$32235 "Waveguide Crossing" sch_x=190 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8252 N$32364 N$32366 N$32237 N$32239 "Waveguide Crossing" sch_x=190 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8253 N$32368 N$32370 N$32241 N$32243 "Waveguide Crossing" sch_x=190 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8254 N$32372 N$32374 N$32245 N$32247 "Waveguide Crossing" sch_x=190 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8255 N$32376 N$32378 N$32249 N$32251 "Waveguide Crossing" sch_x=190 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8256 N$32380 N$32382 N$32253 N$32255 "Waveguide Crossing" sch_x=190 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8257 N$32384 N$32386 N$32257 N$32259 "Waveguide Crossing" sch_x=190 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8258 N$32388 N$32390 N$32261 N$32263 "Waveguide Crossing" sch_x=190 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8259 N$32392 N$32394 N$32265 N$32267 "Waveguide Crossing" sch_x=190 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8260 N$32396 N$32398 N$32269 N$32271 "Waveguide Crossing" sch_x=190 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8261 N$32400 N$32402 N$32273 N$32275 "Waveguide Crossing" sch_x=190 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8262 N$32404 N$32406 N$32277 N$32279 "Waveguide Crossing" sch_x=190 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8263 N$32408 N$32410 N$32281 N$32283 "Waveguide Crossing" sch_x=190 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8264 N$32412 N$32414 N$32285 N$32287 "Waveguide Crossing" sch_x=190 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8265 N$32416 N$32418 N$32289 N$32291 "Waveguide Crossing" sch_x=190 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8266 N$32420 N$32422 N$32293 N$32295 "Waveguide Crossing" sch_x=190 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8267 N$32424 N$32426 N$32297 N$32299 "Waveguide Crossing" sch_x=190 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8268 N$32428 N$32430 N$32301 N$32303 "Waveguide Crossing" sch_x=190 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8269 N$32432 N$32434 N$32305 N$32307 "Waveguide Crossing" sch_x=190 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8270 N$32436 N$32438 N$32309 N$32311 "Waveguide Crossing" sch_x=190 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8271 N$32440 N$32442 N$32313 N$32315 "Waveguide Crossing" sch_x=190 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8272 N$32444 N$34493 N$32317 N$32319 "Waveguide Crossing" sch_x=190 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8273 N$34369 N$32446 N$32321 N$32323 "Waveguide Crossing" sch_x=188 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8274 N$32448 N$32450 N$32325 N$32327 "Waveguide Crossing" sch_x=188 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8275 N$32452 N$32454 N$32329 N$32331 "Waveguide Crossing" sch_x=188 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8276 N$32456 N$32458 N$32333 N$32335 "Waveguide Crossing" sch_x=188 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8277 N$32460 N$32462 N$32337 N$32339 "Waveguide Crossing" sch_x=188 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8278 N$32464 N$32466 N$32341 N$32343 "Waveguide Crossing" sch_x=188 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8279 N$32468 N$32470 N$32345 N$32347 "Waveguide Crossing" sch_x=188 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8280 N$32472 N$32474 N$32349 N$32351 "Waveguide Crossing" sch_x=188 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8281 N$32476 N$32478 N$32353 N$32355 "Waveguide Crossing" sch_x=188 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8282 N$32480 N$32482 N$32357 N$32359 "Waveguide Crossing" sch_x=188 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8283 N$32484 N$32486 N$32361 N$32363 "Waveguide Crossing" sch_x=188 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8284 N$32488 N$32490 N$32365 N$32367 "Waveguide Crossing" sch_x=188 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8285 N$32492 N$32494 N$32369 N$32371 "Waveguide Crossing" sch_x=188 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8286 N$32496 N$32498 N$32373 N$32375 "Waveguide Crossing" sch_x=188 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8287 N$32500 N$32502 N$32377 N$32379 "Waveguide Crossing" sch_x=188 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8288 N$32504 N$32506 N$32381 N$32383 "Waveguide Crossing" sch_x=188 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8289 N$32508 N$32510 N$32385 N$32387 "Waveguide Crossing" sch_x=188 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8290 N$32512 N$32514 N$32389 N$32391 "Waveguide Crossing" sch_x=188 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8291 N$32516 N$32518 N$32393 N$32395 "Waveguide Crossing" sch_x=188 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8292 N$32520 N$32522 N$32397 N$32399 "Waveguide Crossing" sch_x=188 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8293 N$32524 N$32526 N$32401 N$32403 "Waveguide Crossing" sch_x=188 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8294 N$32528 N$32530 N$32405 N$32407 "Waveguide Crossing" sch_x=188 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8295 N$32532 N$32534 N$32409 N$32411 "Waveguide Crossing" sch_x=188 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8296 N$32536 N$32538 N$32413 N$32415 "Waveguide Crossing" sch_x=188 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8297 N$32540 N$32542 N$32417 N$32419 "Waveguide Crossing" sch_x=188 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8298 N$32544 N$32546 N$32421 N$32423 "Waveguide Crossing" sch_x=188 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8299 N$32548 N$32550 N$32425 N$32427 "Waveguide Crossing" sch_x=188 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8300 N$32552 N$32554 N$32429 N$32431 "Waveguide Crossing" sch_x=188 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8301 N$32556 N$32558 N$32433 N$32435 "Waveguide Crossing" sch_x=188 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8302 N$32560 N$32562 N$32437 N$32439 "Waveguide Crossing" sch_x=188 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8303 N$32564 N$34491 N$32441 N$32443 "Waveguide Crossing" sch_x=188 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8304 N$34371 N$32566 N$32445 N$32447 "Waveguide Crossing" sch_x=186 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8305 N$32568 N$32570 N$32449 N$32451 "Waveguide Crossing" sch_x=186 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8306 N$32572 N$32574 N$32453 N$32455 "Waveguide Crossing" sch_x=186 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8307 N$32576 N$32578 N$32457 N$32459 "Waveguide Crossing" sch_x=186 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8308 N$32580 N$32582 N$32461 N$32463 "Waveguide Crossing" sch_x=186 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8309 N$32584 N$32586 N$32465 N$32467 "Waveguide Crossing" sch_x=186 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8310 N$32588 N$32590 N$32469 N$32471 "Waveguide Crossing" sch_x=186 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8311 N$32592 N$32594 N$32473 N$32475 "Waveguide Crossing" sch_x=186 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8312 N$32596 N$32598 N$32477 N$32479 "Waveguide Crossing" sch_x=186 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8313 N$32600 N$32602 N$32481 N$32483 "Waveguide Crossing" sch_x=186 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8314 N$32604 N$32606 N$32485 N$32487 "Waveguide Crossing" sch_x=186 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8315 N$32608 N$32610 N$32489 N$32491 "Waveguide Crossing" sch_x=186 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8316 N$32612 N$32614 N$32493 N$32495 "Waveguide Crossing" sch_x=186 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8317 N$32616 N$32618 N$32497 N$32499 "Waveguide Crossing" sch_x=186 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8318 N$32620 N$32622 N$32501 N$32503 "Waveguide Crossing" sch_x=186 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8319 N$32624 N$32626 N$32505 N$32507 "Waveguide Crossing" sch_x=186 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8320 N$32628 N$32630 N$32509 N$32511 "Waveguide Crossing" sch_x=186 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8321 N$32632 N$32634 N$32513 N$32515 "Waveguide Crossing" sch_x=186 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8322 N$32636 N$32638 N$32517 N$32519 "Waveguide Crossing" sch_x=186 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8323 N$32640 N$32642 N$32521 N$32523 "Waveguide Crossing" sch_x=186 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8324 N$32644 N$32646 N$32525 N$32527 "Waveguide Crossing" sch_x=186 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8325 N$32648 N$32650 N$32529 N$32531 "Waveguide Crossing" sch_x=186 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8326 N$32652 N$32654 N$32533 N$32535 "Waveguide Crossing" sch_x=186 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8327 N$32656 N$32658 N$32537 N$32539 "Waveguide Crossing" sch_x=186 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8328 N$32660 N$32662 N$32541 N$32543 "Waveguide Crossing" sch_x=186 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8329 N$32664 N$32666 N$32545 N$32547 "Waveguide Crossing" sch_x=186 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8330 N$32668 N$32670 N$32549 N$32551 "Waveguide Crossing" sch_x=186 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8331 N$32672 N$32674 N$32553 N$32555 "Waveguide Crossing" sch_x=186 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8332 N$32676 N$32678 N$32557 N$32559 "Waveguide Crossing" sch_x=186 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8333 N$32680 N$34489 N$32561 N$32563 "Waveguide Crossing" sch_x=186 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8334 N$34373 N$32682 N$32565 N$32567 "Waveguide Crossing" sch_x=184 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8335 N$32684 N$32686 N$32569 N$32571 "Waveguide Crossing" sch_x=184 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8336 N$32688 N$32690 N$32573 N$32575 "Waveguide Crossing" sch_x=184 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8337 N$32692 N$32694 N$32577 N$32579 "Waveguide Crossing" sch_x=184 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8338 N$32696 N$32698 N$32581 N$32583 "Waveguide Crossing" sch_x=184 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8339 N$32700 N$32702 N$32585 N$32587 "Waveguide Crossing" sch_x=184 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8340 N$32704 N$32706 N$32589 N$32591 "Waveguide Crossing" sch_x=184 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8341 N$32708 N$32710 N$32593 N$32595 "Waveguide Crossing" sch_x=184 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8342 N$32712 N$32714 N$32597 N$32599 "Waveguide Crossing" sch_x=184 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8343 N$32716 N$32718 N$32601 N$32603 "Waveguide Crossing" sch_x=184 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8344 N$32720 N$32722 N$32605 N$32607 "Waveguide Crossing" sch_x=184 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8345 N$32724 N$32726 N$32609 N$32611 "Waveguide Crossing" sch_x=184 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8346 N$32728 N$32730 N$32613 N$32615 "Waveguide Crossing" sch_x=184 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8347 N$32732 N$32734 N$32617 N$32619 "Waveguide Crossing" sch_x=184 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8348 N$32736 N$32738 N$32621 N$32623 "Waveguide Crossing" sch_x=184 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8349 N$32740 N$32742 N$32625 N$32627 "Waveguide Crossing" sch_x=184 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8350 N$32744 N$32746 N$32629 N$32631 "Waveguide Crossing" sch_x=184 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8351 N$32748 N$32750 N$32633 N$32635 "Waveguide Crossing" sch_x=184 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8352 N$32752 N$32754 N$32637 N$32639 "Waveguide Crossing" sch_x=184 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8353 N$32756 N$32758 N$32641 N$32643 "Waveguide Crossing" sch_x=184 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8354 N$32760 N$32762 N$32645 N$32647 "Waveguide Crossing" sch_x=184 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8355 N$32764 N$32766 N$32649 N$32651 "Waveguide Crossing" sch_x=184 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8356 N$32768 N$32770 N$32653 N$32655 "Waveguide Crossing" sch_x=184 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8357 N$32772 N$32774 N$32657 N$32659 "Waveguide Crossing" sch_x=184 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8358 N$32776 N$32778 N$32661 N$32663 "Waveguide Crossing" sch_x=184 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8359 N$32780 N$32782 N$32665 N$32667 "Waveguide Crossing" sch_x=184 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8360 N$32784 N$32786 N$32669 N$32671 "Waveguide Crossing" sch_x=184 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8361 N$32788 N$32790 N$32673 N$32675 "Waveguide Crossing" sch_x=184 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8362 N$32792 N$34487 N$32677 N$32679 "Waveguide Crossing" sch_x=184 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8363 N$34375 N$32794 N$32681 N$32683 "Waveguide Crossing" sch_x=182 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8364 N$32796 N$32798 N$32685 N$32687 "Waveguide Crossing" sch_x=182 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8365 N$32800 N$32802 N$32689 N$32691 "Waveguide Crossing" sch_x=182 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8366 N$32804 N$32806 N$32693 N$32695 "Waveguide Crossing" sch_x=182 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8367 N$32808 N$32810 N$32697 N$32699 "Waveguide Crossing" sch_x=182 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8368 N$32812 N$32814 N$32701 N$32703 "Waveguide Crossing" sch_x=182 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8369 N$32816 N$32818 N$32705 N$32707 "Waveguide Crossing" sch_x=182 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8370 N$32820 N$32822 N$32709 N$32711 "Waveguide Crossing" sch_x=182 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8371 N$32824 N$32826 N$32713 N$32715 "Waveguide Crossing" sch_x=182 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8372 N$32828 N$32830 N$32717 N$32719 "Waveguide Crossing" sch_x=182 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8373 N$32832 N$32834 N$32721 N$32723 "Waveguide Crossing" sch_x=182 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8374 N$32836 N$32838 N$32725 N$32727 "Waveguide Crossing" sch_x=182 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8375 N$32840 N$32842 N$32729 N$32731 "Waveguide Crossing" sch_x=182 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8376 N$32844 N$32846 N$32733 N$32735 "Waveguide Crossing" sch_x=182 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8377 N$32848 N$32850 N$32737 N$32739 "Waveguide Crossing" sch_x=182 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8378 N$32852 N$32854 N$32741 N$32743 "Waveguide Crossing" sch_x=182 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8379 N$32856 N$32858 N$32745 N$32747 "Waveguide Crossing" sch_x=182 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8380 N$32860 N$32862 N$32749 N$32751 "Waveguide Crossing" sch_x=182 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8381 N$32864 N$32866 N$32753 N$32755 "Waveguide Crossing" sch_x=182 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8382 N$32868 N$32870 N$32757 N$32759 "Waveguide Crossing" sch_x=182 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8383 N$32872 N$32874 N$32761 N$32763 "Waveguide Crossing" sch_x=182 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8384 N$32876 N$32878 N$32765 N$32767 "Waveguide Crossing" sch_x=182 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8385 N$32880 N$32882 N$32769 N$32771 "Waveguide Crossing" sch_x=182 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8386 N$32884 N$32886 N$32773 N$32775 "Waveguide Crossing" sch_x=182 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8387 N$32888 N$32890 N$32777 N$32779 "Waveguide Crossing" sch_x=182 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8388 N$32892 N$32894 N$32781 N$32783 "Waveguide Crossing" sch_x=182 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8389 N$32896 N$32898 N$32785 N$32787 "Waveguide Crossing" sch_x=182 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8390 N$32900 N$34485 N$32789 N$32791 "Waveguide Crossing" sch_x=182 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8391 N$34377 N$32902 N$32793 N$32795 "Waveguide Crossing" sch_x=180 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8392 N$32904 N$32906 N$32797 N$32799 "Waveguide Crossing" sch_x=180 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8393 N$32908 N$32910 N$32801 N$32803 "Waveguide Crossing" sch_x=180 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8394 N$32912 N$32914 N$32805 N$32807 "Waveguide Crossing" sch_x=180 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8395 N$32916 N$32918 N$32809 N$32811 "Waveguide Crossing" sch_x=180 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8396 N$32920 N$32922 N$32813 N$32815 "Waveguide Crossing" sch_x=180 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8397 N$32924 N$32926 N$32817 N$32819 "Waveguide Crossing" sch_x=180 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8398 N$32928 N$32930 N$32821 N$32823 "Waveguide Crossing" sch_x=180 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8399 N$32932 N$32934 N$32825 N$32827 "Waveguide Crossing" sch_x=180 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8400 N$32936 N$32938 N$32829 N$32831 "Waveguide Crossing" sch_x=180 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8401 N$32940 N$32942 N$32833 N$32835 "Waveguide Crossing" sch_x=180 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8402 N$32944 N$32946 N$32837 N$32839 "Waveguide Crossing" sch_x=180 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8403 N$32948 N$32950 N$32841 N$32843 "Waveguide Crossing" sch_x=180 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8404 N$32952 N$32954 N$32845 N$32847 "Waveguide Crossing" sch_x=180 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8405 N$32956 N$32958 N$32849 N$32851 "Waveguide Crossing" sch_x=180 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8406 N$32960 N$32962 N$32853 N$32855 "Waveguide Crossing" sch_x=180 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8407 N$32964 N$32966 N$32857 N$32859 "Waveguide Crossing" sch_x=180 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8408 N$32968 N$32970 N$32861 N$32863 "Waveguide Crossing" sch_x=180 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8409 N$32972 N$32974 N$32865 N$32867 "Waveguide Crossing" sch_x=180 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8410 N$32976 N$32978 N$32869 N$32871 "Waveguide Crossing" sch_x=180 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8411 N$32980 N$32982 N$32873 N$32875 "Waveguide Crossing" sch_x=180 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8412 N$32984 N$32986 N$32877 N$32879 "Waveguide Crossing" sch_x=180 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8413 N$32988 N$32990 N$32881 N$32883 "Waveguide Crossing" sch_x=180 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8414 N$32992 N$32994 N$32885 N$32887 "Waveguide Crossing" sch_x=180 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8415 N$32996 N$32998 N$32889 N$32891 "Waveguide Crossing" sch_x=180 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8416 N$33000 N$33002 N$32893 N$32895 "Waveguide Crossing" sch_x=180 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8417 N$33004 N$34483 N$32897 N$32899 "Waveguide Crossing" sch_x=180 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8418 N$34379 N$33006 N$32901 N$32903 "Waveguide Crossing" sch_x=178 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8419 N$33008 N$33010 N$32905 N$32907 "Waveguide Crossing" sch_x=178 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8420 N$33012 N$33014 N$32909 N$32911 "Waveguide Crossing" sch_x=178 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8421 N$33016 N$33018 N$32913 N$32915 "Waveguide Crossing" sch_x=178 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8422 N$33020 N$33022 N$32917 N$32919 "Waveguide Crossing" sch_x=178 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8423 N$33024 N$33026 N$32921 N$32923 "Waveguide Crossing" sch_x=178 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8424 N$33028 N$33030 N$32925 N$32927 "Waveguide Crossing" sch_x=178 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8425 N$33032 N$33034 N$32929 N$32931 "Waveguide Crossing" sch_x=178 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8426 N$33036 N$33038 N$32933 N$32935 "Waveguide Crossing" sch_x=178 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8427 N$33040 N$33042 N$32937 N$32939 "Waveguide Crossing" sch_x=178 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8428 N$33044 N$33046 N$32941 N$32943 "Waveguide Crossing" sch_x=178 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8429 N$33048 N$33050 N$32945 N$32947 "Waveguide Crossing" sch_x=178 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8430 N$33052 N$33054 N$32949 N$32951 "Waveguide Crossing" sch_x=178 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8431 N$33056 N$33058 N$32953 N$32955 "Waveguide Crossing" sch_x=178 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8432 N$33060 N$33062 N$32957 N$32959 "Waveguide Crossing" sch_x=178 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8433 N$33064 N$33066 N$32961 N$32963 "Waveguide Crossing" sch_x=178 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8434 N$33068 N$33070 N$32965 N$32967 "Waveguide Crossing" sch_x=178 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8435 N$33072 N$33074 N$32969 N$32971 "Waveguide Crossing" sch_x=178 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8436 N$33076 N$33078 N$32973 N$32975 "Waveguide Crossing" sch_x=178 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8437 N$33080 N$33082 N$32977 N$32979 "Waveguide Crossing" sch_x=178 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8438 N$33084 N$33086 N$32981 N$32983 "Waveguide Crossing" sch_x=178 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8439 N$33088 N$33090 N$32985 N$32987 "Waveguide Crossing" sch_x=178 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8440 N$33092 N$33094 N$32989 N$32991 "Waveguide Crossing" sch_x=178 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8441 N$33096 N$33098 N$32993 N$32995 "Waveguide Crossing" sch_x=178 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8442 N$33100 N$33102 N$32997 N$32999 "Waveguide Crossing" sch_x=178 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8443 N$33104 N$34481 N$33001 N$33003 "Waveguide Crossing" sch_x=178 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8444 N$34381 N$33106 N$33005 N$33007 "Waveguide Crossing" sch_x=176 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8445 N$33108 N$33110 N$33009 N$33011 "Waveguide Crossing" sch_x=176 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8446 N$33112 N$33114 N$33013 N$33015 "Waveguide Crossing" sch_x=176 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8447 N$33116 N$33118 N$33017 N$33019 "Waveguide Crossing" sch_x=176 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8448 N$33120 N$33122 N$33021 N$33023 "Waveguide Crossing" sch_x=176 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8449 N$33124 N$33126 N$33025 N$33027 "Waveguide Crossing" sch_x=176 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8450 N$33128 N$33130 N$33029 N$33031 "Waveguide Crossing" sch_x=176 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8451 N$33132 N$33134 N$33033 N$33035 "Waveguide Crossing" sch_x=176 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8452 N$33136 N$33138 N$33037 N$33039 "Waveguide Crossing" sch_x=176 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8453 N$33140 N$33142 N$33041 N$33043 "Waveguide Crossing" sch_x=176 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8454 N$33144 N$33146 N$33045 N$33047 "Waveguide Crossing" sch_x=176 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8455 N$33148 N$33150 N$33049 N$33051 "Waveguide Crossing" sch_x=176 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8456 N$33152 N$33154 N$33053 N$33055 "Waveguide Crossing" sch_x=176 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8457 N$33156 N$33158 N$33057 N$33059 "Waveguide Crossing" sch_x=176 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8458 N$33160 N$33162 N$33061 N$33063 "Waveguide Crossing" sch_x=176 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8459 N$33164 N$33166 N$33065 N$33067 "Waveguide Crossing" sch_x=176 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8460 N$33168 N$33170 N$33069 N$33071 "Waveguide Crossing" sch_x=176 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8461 N$33172 N$33174 N$33073 N$33075 "Waveguide Crossing" sch_x=176 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8462 N$33176 N$33178 N$33077 N$33079 "Waveguide Crossing" sch_x=176 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8463 N$33180 N$33182 N$33081 N$33083 "Waveguide Crossing" sch_x=176 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8464 N$33184 N$33186 N$33085 N$33087 "Waveguide Crossing" sch_x=176 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8465 N$33188 N$33190 N$33089 N$33091 "Waveguide Crossing" sch_x=176 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8466 N$33192 N$33194 N$33093 N$33095 "Waveguide Crossing" sch_x=176 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8467 N$33196 N$33198 N$33097 N$33099 "Waveguide Crossing" sch_x=176 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8468 N$33200 N$34479 N$33101 N$33103 "Waveguide Crossing" sch_x=176 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8469 N$34383 N$33202 N$33105 N$33107 "Waveguide Crossing" sch_x=174 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8470 N$33204 N$33206 N$33109 N$33111 "Waveguide Crossing" sch_x=174 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8471 N$33208 N$33210 N$33113 N$33115 "Waveguide Crossing" sch_x=174 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8472 N$33212 N$33214 N$33117 N$33119 "Waveguide Crossing" sch_x=174 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8473 N$33216 N$33218 N$33121 N$33123 "Waveguide Crossing" sch_x=174 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8474 N$33220 N$33222 N$33125 N$33127 "Waveguide Crossing" sch_x=174 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8475 N$33224 N$33226 N$33129 N$33131 "Waveguide Crossing" sch_x=174 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8476 N$33228 N$33230 N$33133 N$33135 "Waveguide Crossing" sch_x=174 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8477 N$33232 N$33234 N$33137 N$33139 "Waveguide Crossing" sch_x=174 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8478 N$33236 N$33238 N$33141 N$33143 "Waveguide Crossing" sch_x=174 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8479 N$33240 N$33242 N$33145 N$33147 "Waveguide Crossing" sch_x=174 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8480 N$33244 N$33246 N$33149 N$33151 "Waveguide Crossing" sch_x=174 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8481 N$33248 N$33250 N$33153 N$33155 "Waveguide Crossing" sch_x=174 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8482 N$33252 N$33254 N$33157 N$33159 "Waveguide Crossing" sch_x=174 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8483 N$33256 N$33258 N$33161 N$33163 "Waveguide Crossing" sch_x=174 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8484 N$33260 N$33262 N$33165 N$33167 "Waveguide Crossing" sch_x=174 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8485 N$33264 N$33266 N$33169 N$33171 "Waveguide Crossing" sch_x=174 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8486 N$33268 N$33270 N$33173 N$33175 "Waveguide Crossing" sch_x=174 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8487 N$33272 N$33274 N$33177 N$33179 "Waveguide Crossing" sch_x=174 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8488 N$33276 N$33278 N$33181 N$33183 "Waveguide Crossing" sch_x=174 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8489 N$33280 N$33282 N$33185 N$33187 "Waveguide Crossing" sch_x=174 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8490 N$33284 N$33286 N$33189 N$33191 "Waveguide Crossing" sch_x=174 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8491 N$33288 N$33290 N$33193 N$33195 "Waveguide Crossing" sch_x=174 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8492 N$33292 N$34477 N$33197 N$33199 "Waveguide Crossing" sch_x=174 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8493 N$34385 N$33294 N$33201 N$33203 "Waveguide Crossing" sch_x=172 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8494 N$33296 N$33298 N$33205 N$33207 "Waveguide Crossing" sch_x=172 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8495 N$33300 N$33302 N$33209 N$33211 "Waveguide Crossing" sch_x=172 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8496 N$33304 N$33306 N$33213 N$33215 "Waveguide Crossing" sch_x=172 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8497 N$33308 N$33310 N$33217 N$33219 "Waveguide Crossing" sch_x=172 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8498 N$33312 N$33314 N$33221 N$33223 "Waveguide Crossing" sch_x=172 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8499 N$33316 N$33318 N$33225 N$33227 "Waveguide Crossing" sch_x=172 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8500 N$33320 N$33322 N$33229 N$33231 "Waveguide Crossing" sch_x=172 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8501 N$33324 N$33326 N$33233 N$33235 "Waveguide Crossing" sch_x=172 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8502 N$33328 N$33330 N$33237 N$33239 "Waveguide Crossing" sch_x=172 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8503 N$33332 N$33334 N$33241 N$33243 "Waveguide Crossing" sch_x=172 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8504 N$33336 N$33338 N$33245 N$33247 "Waveguide Crossing" sch_x=172 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8505 N$33340 N$33342 N$33249 N$33251 "Waveguide Crossing" sch_x=172 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8506 N$33344 N$33346 N$33253 N$33255 "Waveguide Crossing" sch_x=172 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8507 N$33348 N$33350 N$33257 N$33259 "Waveguide Crossing" sch_x=172 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8508 N$33352 N$33354 N$33261 N$33263 "Waveguide Crossing" sch_x=172 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8509 N$33356 N$33358 N$33265 N$33267 "Waveguide Crossing" sch_x=172 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8510 N$33360 N$33362 N$33269 N$33271 "Waveguide Crossing" sch_x=172 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8511 N$33364 N$33366 N$33273 N$33275 "Waveguide Crossing" sch_x=172 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8512 N$33368 N$33370 N$33277 N$33279 "Waveguide Crossing" sch_x=172 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8513 N$33372 N$33374 N$33281 N$33283 "Waveguide Crossing" sch_x=172 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8514 N$33376 N$33378 N$33285 N$33287 "Waveguide Crossing" sch_x=172 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8515 N$33380 N$34475 N$33289 N$33291 "Waveguide Crossing" sch_x=172 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8516 N$34387 N$33382 N$33293 N$33295 "Waveguide Crossing" sch_x=170 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8517 N$33384 N$33386 N$33297 N$33299 "Waveguide Crossing" sch_x=170 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8518 N$33388 N$33390 N$33301 N$33303 "Waveguide Crossing" sch_x=170 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8519 N$33392 N$33394 N$33305 N$33307 "Waveguide Crossing" sch_x=170 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8520 N$33396 N$33398 N$33309 N$33311 "Waveguide Crossing" sch_x=170 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8521 N$33400 N$33402 N$33313 N$33315 "Waveguide Crossing" sch_x=170 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8522 N$33404 N$33406 N$33317 N$33319 "Waveguide Crossing" sch_x=170 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8523 N$33408 N$33410 N$33321 N$33323 "Waveguide Crossing" sch_x=170 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8524 N$33412 N$33414 N$33325 N$33327 "Waveguide Crossing" sch_x=170 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8525 N$33416 N$33418 N$33329 N$33331 "Waveguide Crossing" sch_x=170 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8526 N$33420 N$33422 N$33333 N$33335 "Waveguide Crossing" sch_x=170 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8527 N$33424 N$33426 N$33337 N$33339 "Waveguide Crossing" sch_x=170 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8528 N$33428 N$33430 N$33341 N$33343 "Waveguide Crossing" sch_x=170 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8529 N$33432 N$33434 N$33345 N$33347 "Waveguide Crossing" sch_x=170 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8530 N$33436 N$33438 N$33349 N$33351 "Waveguide Crossing" sch_x=170 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8531 N$33440 N$33442 N$33353 N$33355 "Waveguide Crossing" sch_x=170 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8532 N$33444 N$33446 N$33357 N$33359 "Waveguide Crossing" sch_x=170 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8533 N$33448 N$33450 N$33361 N$33363 "Waveguide Crossing" sch_x=170 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8534 N$33452 N$33454 N$33365 N$33367 "Waveguide Crossing" sch_x=170 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8535 N$33456 N$33458 N$33369 N$33371 "Waveguide Crossing" sch_x=170 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8536 N$33460 N$33462 N$33373 N$33375 "Waveguide Crossing" sch_x=170 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8537 N$33464 N$34473 N$33377 N$33379 "Waveguide Crossing" sch_x=170 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8538 N$34389 N$33466 N$33381 N$33383 "Waveguide Crossing" sch_x=168 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8539 N$33468 N$33470 N$33385 N$33387 "Waveguide Crossing" sch_x=168 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8540 N$33472 N$33474 N$33389 N$33391 "Waveguide Crossing" sch_x=168 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8541 N$33476 N$33478 N$33393 N$33395 "Waveguide Crossing" sch_x=168 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8542 N$33480 N$33482 N$33397 N$33399 "Waveguide Crossing" sch_x=168 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8543 N$33484 N$33486 N$33401 N$33403 "Waveguide Crossing" sch_x=168 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8544 N$33488 N$33490 N$33405 N$33407 "Waveguide Crossing" sch_x=168 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8545 N$33492 N$33494 N$33409 N$33411 "Waveguide Crossing" sch_x=168 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8546 N$33496 N$33498 N$33413 N$33415 "Waveguide Crossing" sch_x=168 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8547 N$33500 N$33502 N$33417 N$33419 "Waveguide Crossing" sch_x=168 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8548 N$33504 N$33506 N$33421 N$33423 "Waveguide Crossing" sch_x=168 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8549 N$33508 N$33510 N$33425 N$33427 "Waveguide Crossing" sch_x=168 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8550 N$33512 N$33514 N$33429 N$33431 "Waveguide Crossing" sch_x=168 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8551 N$33516 N$33518 N$33433 N$33435 "Waveguide Crossing" sch_x=168 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8552 N$33520 N$33522 N$33437 N$33439 "Waveguide Crossing" sch_x=168 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8553 N$33524 N$33526 N$33441 N$33443 "Waveguide Crossing" sch_x=168 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8554 N$33528 N$33530 N$33445 N$33447 "Waveguide Crossing" sch_x=168 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8555 N$33532 N$33534 N$33449 N$33451 "Waveguide Crossing" sch_x=168 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8556 N$33536 N$33538 N$33453 N$33455 "Waveguide Crossing" sch_x=168 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8557 N$33540 N$33542 N$33457 N$33459 "Waveguide Crossing" sch_x=168 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8558 N$33544 N$34471 N$33461 N$33463 "Waveguide Crossing" sch_x=168 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8559 N$34391 N$33546 N$33465 N$33467 "Waveguide Crossing" sch_x=166 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8560 N$33548 N$33550 N$33469 N$33471 "Waveguide Crossing" sch_x=166 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8561 N$33552 N$33554 N$33473 N$33475 "Waveguide Crossing" sch_x=166 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8562 N$33556 N$33558 N$33477 N$33479 "Waveguide Crossing" sch_x=166 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8563 N$33560 N$33562 N$33481 N$33483 "Waveguide Crossing" sch_x=166 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8564 N$33564 N$33566 N$33485 N$33487 "Waveguide Crossing" sch_x=166 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8565 N$33568 N$33570 N$33489 N$33491 "Waveguide Crossing" sch_x=166 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8566 N$33572 N$33574 N$33493 N$33495 "Waveguide Crossing" sch_x=166 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8567 N$33576 N$33578 N$33497 N$33499 "Waveguide Crossing" sch_x=166 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8568 N$33580 N$33582 N$33501 N$33503 "Waveguide Crossing" sch_x=166 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8569 N$33584 N$33586 N$33505 N$33507 "Waveguide Crossing" sch_x=166 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8570 N$33588 N$33590 N$33509 N$33511 "Waveguide Crossing" sch_x=166 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8571 N$33592 N$33594 N$33513 N$33515 "Waveguide Crossing" sch_x=166 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8572 N$33596 N$33598 N$33517 N$33519 "Waveguide Crossing" sch_x=166 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8573 N$33600 N$33602 N$33521 N$33523 "Waveguide Crossing" sch_x=166 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8574 N$33604 N$33606 N$33525 N$33527 "Waveguide Crossing" sch_x=166 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8575 N$33608 N$33610 N$33529 N$33531 "Waveguide Crossing" sch_x=166 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8576 N$33612 N$33614 N$33533 N$33535 "Waveguide Crossing" sch_x=166 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8577 N$33616 N$33618 N$33537 N$33539 "Waveguide Crossing" sch_x=166 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8578 N$33620 N$34469 N$33541 N$33543 "Waveguide Crossing" sch_x=166 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8579 N$34393 N$33622 N$33545 N$33547 "Waveguide Crossing" sch_x=164 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8580 N$33624 N$33626 N$33549 N$33551 "Waveguide Crossing" sch_x=164 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8581 N$33628 N$33630 N$33553 N$33555 "Waveguide Crossing" sch_x=164 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8582 N$33632 N$33634 N$33557 N$33559 "Waveguide Crossing" sch_x=164 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8583 N$33636 N$33638 N$33561 N$33563 "Waveguide Crossing" sch_x=164 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8584 N$33640 N$33642 N$33565 N$33567 "Waveguide Crossing" sch_x=164 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8585 N$33644 N$33646 N$33569 N$33571 "Waveguide Crossing" sch_x=164 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8586 N$33648 N$33650 N$33573 N$33575 "Waveguide Crossing" sch_x=164 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8587 N$33652 N$33654 N$33577 N$33579 "Waveguide Crossing" sch_x=164 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8588 N$33656 N$33658 N$33581 N$33583 "Waveguide Crossing" sch_x=164 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8589 N$33660 N$33662 N$33585 N$33587 "Waveguide Crossing" sch_x=164 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8590 N$33664 N$33666 N$33589 N$33591 "Waveguide Crossing" sch_x=164 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8591 N$33668 N$33670 N$33593 N$33595 "Waveguide Crossing" sch_x=164 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8592 N$33672 N$33674 N$33597 N$33599 "Waveguide Crossing" sch_x=164 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8593 N$33676 N$33678 N$33601 N$33603 "Waveguide Crossing" sch_x=164 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8594 N$33680 N$33682 N$33605 N$33607 "Waveguide Crossing" sch_x=164 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8595 N$33684 N$33686 N$33609 N$33611 "Waveguide Crossing" sch_x=164 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8596 N$33688 N$33690 N$33613 N$33615 "Waveguide Crossing" sch_x=164 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8597 N$33692 N$34467 N$33617 N$33619 "Waveguide Crossing" sch_x=164 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8598 N$34395 N$33694 N$33621 N$33623 "Waveguide Crossing" sch_x=162 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8599 N$33696 N$33698 N$33625 N$33627 "Waveguide Crossing" sch_x=162 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8600 N$33700 N$33702 N$33629 N$33631 "Waveguide Crossing" sch_x=162 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8601 N$33704 N$33706 N$33633 N$33635 "Waveguide Crossing" sch_x=162 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8602 N$33708 N$33710 N$33637 N$33639 "Waveguide Crossing" sch_x=162 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8603 N$33712 N$33714 N$33641 N$33643 "Waveguide Crossing" sch_x=162 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8604 N$33716 N$33718 N$33645 N$33647 "Waveguide Crossing" sch_x=162 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8605 N$33720 N$33722 N$33649 N$33651 "Waveguide Crossing" sch_x=162 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8606 N$33724 N$33726 N$33653 N$33655 "Waveguide Crossing" sch_x=162 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8607 N$33728 N$33730 N$33657 N$33659 "Waveguide Crossing" sch_x=162 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8608 N$33732 N$33734 N$33661 N$33663 "Waveguide Crossing" sch_x=162 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8609 N$33736 N$33738 N$33665 N$33667 "Waveguide Crossing" sch_x=162 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8610 N$33740 N$33742 N$33669 N$33671 "Waveguide Crossing" sch_x=162 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8611 N$33744 N$33746 N$33673 N$33675 "Waveguide Crossing" sch_x=162 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8612 N$33748 N$33750 N$33677 N$33679 "Waveguide Crossing" sch_x=162 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8613 N$33752 N$33754 N$33681 N$33683 "Waveguide Crossing" sch_x=162 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8614 N$33756 N$33758 N$33685 N$33687 "Waveguide Crossing" sch_x=162 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8615 N$33760 N$34465 N$33689 N$33691 "Waveguide Crossing" sch_x=162 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8616 N$34397 N$33762 N$33693 N$33695 "Waveguide Crossing" sch_x=160 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8617 N$33764 N$33766 N$33697 N$33699 "Waveguide Crossing" sch_x=160 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8618 N$33768 N$33770 N$33701 N$33703 "Waveguide Crossing" sch_x=160 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8619 N$33772 N$33774 N$33705 N$33707 "Waveguide Crossing" sch_x=160 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8620 N$33776 N$33778 N$33709 N$33711 "Waveguide Crossing" sch_x=160 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8621 N$33780 N$33782 N$33713 N$33715 "Waveguide Crossing" sch_x=160 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8622 N$33784 N$33786 N$33717 N$33719 "Waveguide Crossing" sch_x=160 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8623 N$33788 N$33790 N$33721 N$33723 "Waveguide Crossing" sch_x=160 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8624 N$33792 N$33794 N$33725 N$33727 "Waveguide Crossing" sch_x=160 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8625 N$33796 N$33798 N$33729 N$33731 "Waveguide Crossing" sch_x=160 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8626 N$33800 N$33802 N$33733 N$33735 "Waveguide Crossing" sch_x=160 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8627 N$33804 N$33806 N$33737 N$33739 "Waveguide Crossing" sch_x=160 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8628 N$33808 N$33810 N$33741 N$33743 "Waveguide Crossing" sch_x=160 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8629 N$33812 N$33814 N$33745 N$33747 "Waveguide Crossing" sch_x=160 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8630 N$33816 N$33818 N$33749 N$33751 "Waveguide Crossing" sch_x=160 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8631 N$33820 N$33822 N$33753 N$33755 "Waveguide Crossing" sch_x=160 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8632 N$33824 N$34463 N$33757 N$33759 "Waveguide Crossing" sch_x=160 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8633 N$34399 N$33826 N$33761 N$33763 "Waveguide Crossing" sch_x=158 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8634 N$33828 N$33830 N$33765 N$33767 "Waveguide Crossing" sch_x=158 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8635 N$33832 N$33834 N$33769 N$33771 "Waveguide Crossing" sch_x=158 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8636 N$33836 N$33838 N$33773 N$33775 "Waveguide Crossing" sch_x=158 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8637 N$33840 N$33842 N$33777 N$33779 "Waveguide Crossing" sch_x=158 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8638 N$33844 N$33846 N$33781 N$33783 "Waveguide Crossing" sch_x=158 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8639 N$33848 N$33850 N$33785 N$33787 "Waveguide Crossing" sch_x=158 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8640 N$33852 N$33854 N$33789 N$33791 "Waveguide Crossing" sch_x=158 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8641 N$33856 N$33858 N$33793 N$33795 "Waveguide Crossing" sch_x=158 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8642 N$33860 N$33862 N$33797 N$33799 "Waveguide Crossing" sch_x=158 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8643 N$33864 N$33866 N$33801 N$33803 "Waveguide Crossing" sch_x=158 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8644 N$33868 N$33870 N$33805 N$33807 "Waveguide Crossing" sch_x=158 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8645 N$33872 N$33874 N$33809 N$33811 "Waveguide Crossing" sch_x=158 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8646 N$33876 N$33878 N$33813 N$33815 "Waveguide Crossing" sch_x=158 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8647 N$33880 N$33882 N$33817 N$33819 "Waveguide Crossing" sch_x=158 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8648 N$33884 N$34461 N$33821 N$33823 "Waveguide Crossing" sch_x=158 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8649 N$34401 N$33886 N$33825 N$33827 "Waveguide Crossing" sch_x=156 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8650 N$33888 N$33890 N$33829 N$33831 "Waveguide Crossing" sch_x=156 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8651 N$33892 N$33894 N$33833 N$33835 "Waveguide Crossing" sch_x=156 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8652 N$33896 N$33898 N$33837 N$33839 "Waveguide Crossing" sch_x=156 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8653 N$33900 N$33902 N$33841 N$33843 "Waveguide Crossing" sch_x=156 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8654 N$33904 N$33906 N$33845 N$33847 "Waveguide Crossing" sch_x=156 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8655 N$33908 N$33910 N$33849 N$33851 "Waveguide Crossing" sch_x=156 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8656 N$33912 N$33914 N$33853 N$33855 "Waveguide Crossing" sch_x=156 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8657 N$33916 N$33918 N$33857 N$33859 "Waveguide Crossing" sch_x=156 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8658 N$33920 N$33922 N$33861 N$33863 "Waveguide Crossing" sch_x=156 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8659 N$33924 N$33926 N$33865 N$33867 "Waveguide Crossing" sch_x=156 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8660 N$33928 N$33930 N$33869 N$33871 "Waveguide Crossing" sch_x=156 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8661 N$33932 N$33934 N$33873 N$33875 "Waveguide Crossing" sch_x=156 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8662 N$33936 N$33938 N$33877 N$33879 "Waveguide Crossing" sch_x=156 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8663 N$33940 N$34459 N$33881 N$33883 "Waveguide Crossing" sch_x=156 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8664 N$34403 N$33942 N$33885 N$33887 "Waveguide Crossing" sch_x=154 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8665 N$33944 N$33946 N$33889 N$33891 "Waveguide Crossing" sch_x=154 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8666 N$33948 N$33950 N$33893 N$33895 "Waveguide Crossing" sch_x=154 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8667 N$33952 N$33954 N$33897 N$33899 "Waveguide Crossing" sch_x=154 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8668 N$33956 N$33958 N$33901 N$33903 "Waveguide Crossing" sch_x=154 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8669 N$33960 N$33962 N$33905 N$33907 "Waveguide Crossing" sch_x=154 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8670 N$33964 N$33966 N$33909 N$33911 "Waveguide Crossing" sch_x=154 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8671 N$33968 N$33970 N$33913 N$33915 "Waveguide Crossing" sch_x=154 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8672 N$33972 N$33974 N$33917 N$33919 "Waveguide Crossing" sch_x=154 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8673 N$33976 N$33978 N$33921 N$33923 "Waveguide Crossing" sch_x=154 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8674 N$33980 N$33982 N$33925 N$33927 "Waveguide Crossing" sch_x=154 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8675 N$33984 N$33986 N$33929 N$33931 "Waveguide Crossing" sch_x=154 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8676 N$33988 N$33990 N$33933 N$33935 "Waveguide Crossing" sch_x=154 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8677 N$33992 N$34457 N$33937 N$33939 "Waveguide Crossing" sch_x=154 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8678 N$34405 N$33994 N$33941 N$33943 "Waveguide Crossing" sch_x=152 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8679 N$33996 N$33998 N$33945 N$33947 "Waveguide Crossing" sch_x=152 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8680 N$34000 N$34002 N$33949 N$33951 "Waveguide Crossing" sch_x=152 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8681 N$34004 N$34006 N$33953 N$33955 "Waveguide Crossing" sch_x=152 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8682 N$34008 N$34010 N$33957 N$33959 "Waveguide Crossing" sch_x=152 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8683 N$34012 N$34014 N$33961 N$33963 "Waveguide Crossing" sch_x=152 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8684 N$34016 N$34018 N$33965 N$33967 "Waveguide Crossing" sch_x=152 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8685 N$34020 N$34022 N$33969 N$33971 "Waveguide Crossing" sch_x=152 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8686 N$34024 N$34026 N$33973 N$33975 "Waveguide Crossing" sch_x=152 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8687 N$34028 N$34030 N$33977 N$33979 "Waveguide Crossing" sch_x=152 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8688 N$34032 N$34034 N$33981 N$33983 "Waveguide Crossing" sch_x=152 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8689 N$34036 N$34038 N$33985 N$33987 "Waveguide Crossing" sch_x=152 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8690 N$34040 N$34455 N$33989 N$33991 "Waveguide Crossing" sch_x=152 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8691 N$34407 N$34042 N$33993 N$33995 "Waveguide Crossing" sch_x=150 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8692 N$34044 N$34046 N$33997 N$33999 "Waveguide Crossing" sch_x=150 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8693 N$34048 N$34050 N$34001 N$34003 "Waveguide Crossing" sch_x=150 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8694 N$34052 N$34054 N$34005 N$34007 "Waveguide Crossing" sch_x=150 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8695 N$34056 N$34058 N$34009 N$34011 "Waveguide Crossing" sch_x=150 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8696 N$34060 N$34062 N$34013 N$34015 "Waveguide Crossing" sch_x=150 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8697 N$34064 N$34066 N$34017 N$34019 "Waveguide Crossing" sch_x=150 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8698 N$34068 N$34070 N$34021 N$34023 "Waveguide Crossing" sch_x=150 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8699 N$34072 N$34074 N$34025 N$34027 "Waveguide Crossing" sch_x=150 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8700 N$34076 N$34078 N$34029 N$34031 "Waveguide Crossing" sch_x=150 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8701 N$34080 N$34082 N$34033 N$34035 "Waveguide Crossing" sch_x=150 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8702 N$34084 N$34453 N$34037 N$34039 "Waveguide Crossing" sch_x=150 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8703 N$34409 N$34086 N$34041 N$34043 "Waveguide Crossing" sch_x=148 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8704 N$34088 N$34090 N$34045 N$34047 "Waveguide Crossing" sch_x=148 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8705 N$34092 N$34094 N$34049 N$34051 "Waveguide Crossing" sch_x=148 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8706 N$34096 N$34098 N$34053 N$34055 "Waveguide Crossing" sch_x=148 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8707 N$34100 N$34102 N$34057 N$34059 "Waveguide Crossing" sch_x=148 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8708 N$34104 N$34106 N$34061 N$34063 "Waveguide Crossing" sch_x=148 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8709 N$34108 N$34110 N$34065 N$34067 "Waveguide Crossing" sch_x=148 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8710 N$34112 N$34114 N$34069 N$34071 "Waveguide Crossing" sch_x=148 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8711 N$34116 N$34118 N$34073 N$34075 "Waveguide Crossing" sch_x=148 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8712 N$34120 N$34122 N$34077 N$34079 "Waveguide Crossing" sch_x=148 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8713 N$34124 N$34451 N$34081 N$34083 "Waveguide Crossing" sch_x=148 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8714 N$34411 N$34126 N$34085 N$34087 "Waveguide Crossing" sch_x=146 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8715 N$34128 N$34130 N$34089 N$34091 "Waveguide Crossing" sch_x=146 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8716 N$34132 N$34134 N$34093 N$34095 "Waveguide Crossing" sch_x=146 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8717 N$34136 N$34138 N$34097 N$34099 "Waveguide Crossing" sch_x=146 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8718 N$34140 N$34142 N$34101 N$34103 "Waveguide Crossing" sch_x=146 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8719 N$34144 N$34146 N$34105 N$34107 "Waveguide Crossing" sch_x=146 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8720 N$34148 N$34150 N$34109 N$34111 "Waveguide Crossing" sch_x=146 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8721 N$34152 N$34154 N$34113 N$34115 "Waveguide Crossing" sch_x=146 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8722 N$34156 N$34158 N$34117 N$34119 "Waveguide Crossing" sch_x=146 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8723 N$34160 N$34449 N$34121 N$34123 "Waveguide Crossing" sch_x=146 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8724 N$34413 N$34162 N$34125 N$34127 "Waveguide Crossing" sch_x=144 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8725 N$34164 N$34166 N$34129 N$34131 "Waveguide Crossing" sch_x=144 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8726 N$34168 N$34170 N$34133 N$34135 "Waveguide Crossing" sch_x=144 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8727 N$34172 N$34174 N$34137 N$34139 "Waveguide Crossing" sch_x=144 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8728 N$34176 N$34178 N$34141 N$34143 "Waveguide Crossing" sch_x=144 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8729 N$34180 N$34182 N$34145 N$34147 "Waveguide Crossing" sch_x=144 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8730 N$34184 N$34186 N$34149 N$34151 "Waveguide Crossing" sch_x=144 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8731 N$34188 N$34190 N$34153 N$34155 "Waveguide Crossing" sch_x=144 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8732 N$34192 N$34447 N$34157 N$34159 "Waveguide Crossing" sch_x=144 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8733 N$34415 N$34194 N$34161 N$34163 "Waveguide Crossing" sch_x=142 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8734 N$34196 N$34198 N$34165 N$34167 "Waveguide Crossing" sch_x=142 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8735 N$34200 N$34202 N$34169 N$34171 "Waveguide Crossing" sch_x=142 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8736 N$34204 N$34206 N$34173 N$34175 "Waveguide Crossing" sch_x=142 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8737 N$34208 N$34210 N$34177 N$34179 "Waveguide Crossing" sch_x=142 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8738 N$34212 N$34214 N$34181 N$34183 "Waveguide Crossing" sch_x=142 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8739 N$34216 N$34218 N$34185 N$34187 "Waveguide Crossing" sch_x=142 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8740 N$34220 N$34445 N$34189 N$34191 "Waveguide Crossing" sch_x=142 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8741 N$34417 N$34222 N$34193 N$34195 "Waveguide Crossing" sch_x=140 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8742 N$34224 N$34226 N$34197 N$34199 "Waveguide Crossing" sch_x=140 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8743 N$34228 N$34230 N$34201 N$34203 "Waveguide Crossing" sch_x=140 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8744 N$34232 N$34234 N$34205 N$34207 "Waveguide Crossing" sch_x=140 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8745 N$34236 N$34238 N$34209 N$34211 "Waveguide Crossing" sch_x=140 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8746 N$34240 N$34242 N$34213 N$34215 "Waveguide Crossing" sch_x=140 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8747 N$34244 N$34443 N$34217 N$34219 "Waveguide Crossing" sch_x=140 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8748 N$34419 N$34246 N$34221 N$34223 "Waveguide Crossing" sch_x=138 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8749 N$34248 N$34250 N$34225 N$34227 "Waveguide Crossing" sch_x=138 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8750 N$34252 N$34254 N$34229 N$34231 "Waveguide Crossing" sch_x=138 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8751 N$34256 N$34258 N$34233 N$34235 "Waveguide Crossing" sch_x=138 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8752 N$34260 N$34262 N$34237 N$34239 "Waveguide Crossing" sch_x=138 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8753 N$34264 N$34441 N$34241 N$34243 "Waveguide Crossing" sch_x=138 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8754 N$34421 N$34266 N$34245 N$34247 "Waveguide Crossing" sch_x=136 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8755 N$34268 N$34270 N$34249 N$34251 "Waveguide Crossing" sch_x=136 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8756 N$34272 N$34274 N$34253 N$34255 "Waveguide Crossing" sch_x=136 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8757 N$34276 N$34278 N$34257 N$34259 "Waveguide Crossing" sch_x=136 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8758 N$34280 N$34439 N$34261 N$34263 "Waveguide Crossing" sch_x=136 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8759 N$34423 N$34282 N$34265 N$34267 "Waveguide Crossing" sch_x=134 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8760 N$34284 N$34286 N$34269 N$34271 "Waveguide Crossing" sch_x=134 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8761 N$34288 N$34290 N$34273 N$34275 "Waveguide Crossing" sch_x=134 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8762 N$34292 N$34437 N$34277 N$34279 "Waveguide Crossing" sch_x=134 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8763 N$34425 N$34294 N$34281 N$34283 "Waveguide Crossing" sch_x=132 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8764 N$34296 N$34298 N$34285 N$34287 "Waveguide Crossing" sch_x=132 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8765 N$34300 N$34435 N$34289 N$34291 "Waveguide Crossing" sch_x=132 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8766 N$34427 N$34302 N$34293 N$34295 "Waveguide Crossing" sch_x=130 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8767 N$34304 N$34433 N$34297 N$34299 "Waveguide Crossing" sch_x=130 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C8768 N$34429 N$34431 N$34301 N$34303 "Waveguide Crossing" sch_x=128 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6689 N$34557 N$26242 N$34945 N$34946 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6690 N$26244 N$26246 N$34947 N$34948 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6691 N$26248 N$26250 N$34949 N$34950 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6692 N$26252 N$26254 N$34951 N$34952 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6693 N$26256 N$26258 N$34953 N$34954 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6694 N$26260 N$26262 N$34955 N$34956 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6695 N$26264 N$26266 N$34957 N$34958 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6696 N$26268 N$26270 N$34959 N$34960 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6697 N$26272 N$26274 N$34961 N$34962 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6698 N$26276 N$26278 N$34963 N$34964 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6699 N$26280 N$26282 N$34965 N$34966 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6700 N$26284 N$26286 N$34967 N$34968 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6701 N$26288 N$26290 N$34969 N$34970 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6702 N$26292 N$26294 N$34971 N$34972 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6703 N$26296 N$26298 N$34973 N$34974 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6704 N$26300 N$26302 N$34975 N$34976 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6705 N$26304 N$26306 N$34977 N$34978 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6706 N$26308 N$26310 N$34979 N$34980 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6707 N$26312 N$26314 N$34981 N$34982 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6708 N$26316 N$26318 N$34983 N$34984 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6709 N$26320 N$26322 N$34985 N$34986 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6710 N$26324 N$26326 N$34987 N$34988 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6711 N$26328 N$26330 N$34989 N$34990 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6712 N$26332 N$26334 N$34991 N$34992 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6713 N$26336 N$26338 N$34993 N$34994 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6714 N$26340 N$26342 N$34995 N$34996 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6715 N$26344 N$26346 N$34997 N$34998 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6716 N$26348 N$26350 N$34999 N$35000 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6717 N$26352 N$26354 N$35001 N$35002 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6718 N$26356 N$26358 N$35003 N$35004 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6719 N$26360 N$26362 N$35005 N$35006 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6720 N$26364 N$26366 N$35007 N$35008 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6721 N$26368 N$26370 N$35009 N$35010 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6722 N$26372 N$26374 N$35011 N$35012 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6723 N$26376 N$26378 N$35013 N$35014 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6724 N$26380 N$26382 N$35015 N$35016 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6725 N$26384 N$26386 N$35017 N$35018 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6726 N$26388 N$26390 N$35019 N$35020 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6727 N$26392 N$26394 N$35021 N$35022 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6728 N$26396 N$26398 N$35023 N$35024 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6729 N$26400 N$26402 N$35025 N$35026 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6730 N$26404 N$26406 N$35027 N$35028 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6731 N$26408 N$26410 N$35029 N$35030 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6732 N$26412 N$26414 N$35031 N$35032 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6733 N$26416 N$26418 N$35033 N$35034 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6734 N$26420 N$26422 N$35035 N$35036 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6735 N$26424 N$26426 N$35037 N$35038 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6736 N$26428 N$26430 N$35039 N$35040 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6737 N$26432 N$26434 N$35041 N$35042 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6738 N$26436 N$26438 N$35043 N$35044 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6739 N$26440 N$26442 N$35045 N$35046 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6740 N$26444 N$26446 N$35047 N$35048 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6741 N$26448 N$26450 N$35049 N$35050 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6742 N$26452 N$26454 N$35051 N$35052 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6743 N$26456 N$26458 N$35053 N$35054 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6744 N$26460 N$26462 N$35055 N$35056 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6745 N$26464 N$26466 N$35057 N$35058 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6746 N$26468 N$26470 N$35059 N$35060 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6747 N$26472 N$26474 N$35061 N$35062 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6748 N$26476 N$26478 N$35063 N$35064 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6749 N$26480 N$26482 N$35065 N$35066 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6750 N$26484 N$26486 N$35067 N$35068 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6751 N$26488 N$26490 N$35069 N$35070 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6752 N$26492 N$34559 N$35071 N$35072 BDC_switch_ideal library="Design kits/capstone" sch_x=254 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1 N$1 N$2 "Straight Waveguide" sch_x=-4 sch_y=63.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2 N$3 N$4 "Straight Waveguide" sch_x=-5 sch_y=62.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3 N$5 N$6 "Straight Waveguide" sch_x=-5 sch_y=61.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4 N$7 N$8 "Straight Waveguide" sch_x=-3 sch_y=62.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5 N$9 N$10 "Straight Waveguide" sch_x=-3 sch_y=61.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6 N$11 N$12 "Straight Waveguide" sch_x=-4 sch_y=60.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7 N$13 N$14 "Straight Waveguide" sch_x=0 sch_y=63.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8 N$15 N$16 "Straight Waveguide" sch_x=-1 sch_y=63.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9 N$17 N$18 "Straight Waveguide" sch_x=-1 sch_y=62.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10 N$19 N$20 "Straight Waveguide" sch_x=1 sch_y=62.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11 N$21 N$22 "Straight Waveguide" sch_x=1 sch_y=63.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12 N$23 N$24 "Straight Waveguide" sch_x=0 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13 N$25 N$26 "Straight Waveguide" sch_x=0 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14 N$27 N$28 "Straight Waveguide" sch_x=-1 sch_y=61.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15 N$29 N$30 "Straight Waveguide" sch_x=-1 sch_y=60.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16 N$31 N$32 "Straight Waveguide" sch_x=1 sch_y=60.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17 N$33 N$34 "Straight Waveguide" sch_x=1 sch_y=61.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W18 N$35 N$36 "Straight Waveguide" sch_x=0 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W19 N$37 N$38 "Straight Waveguide" sch_x=4 sch_y=63.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W20 N$39 N$40 "Straight Waveguide" sch_x=3 sch_y=62.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W21 N$41 N$42 "Straight Waveguide" sch_x=3 sch_y=61.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W22 N$43 N$44 "Straight Waveguide" sch_x=5 sch_y=61.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W23 N$45 N$46 "Straight Waveguide" sch_x=5 sch_y=62.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W24 N$47 N$48 "Straight Waveguide" sch_x=4 sch_y=60.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W25 N$49 N$50 "Straight Waveguide" sch_x=-4 sch_y=59.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W26 N$51 N$52 "Straight Waveguide" sch_x=-5 sch_y=58.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W27 N$53 N$54 "Straight Waveguide" sch_x=-5 sch_y=57.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W28 N$55 N$56 "Straight Waveguide" sch_x=-3 sch_y=58.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W29 N$57 N$58 "Straight Waveguide" sch_x=-3 sch_y=57.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W30 N$59 N$60 "Straight Waveguide" sch_x=-4 sch_y=56.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W31 N$61 N$62 "Straight Waveguide" sch_x=0 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W32 N$63 N$64 "Straight Waveguide" sch_x=-1 sch_y=59.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W33 N$65 N$66 "Straight Waveguide" sch_x=-1 sch_y=58.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W34 N$67 N$68 "Straight Waveguide" sch_x=1 sch_y=58.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W35 N$69 N$70 "Straight Waveguide" sch_x=1 sch_y=59.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W36 N$71 N$72 "Straight Waveguide" sch_x=0 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W37 N$73 N$74 "Straight Waveguide" sch_x=0 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W38 N$75 N$76 "Straight Waveguide" sch_x=-1 sch_y=57.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W39 N$77 N$78 "Straight Waveguide" sch_x=-1 sch_y=56.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W40 N$79 N$80 "Straight Waveguide" sch_x=1 sch_y=56.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W41 N$81 N$82 "Straight Waveguide" sch_x=1 sch_y=57.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W42 N$83 N$84 "Straight Waveguide" sch_x=0 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W43 N$85 N$86 "Straight Waveguide" sch_x=4 sch_y=59.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W44 N$87 N$88 "Straight Waveguide" sch_x=3 sch_y=58.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W45 N$89 N$90 "Straight Waveguide" sch_x=3 sch_y=57.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W46 N$91 N$92 "Straight Waveguide" sch_x=5 sch_y=57.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W47 N$93 N$94 "Straight Waveguide" sch_x=5 sch_y=58.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W48 N$95 N$96 "Straight Waveguide" sch_x=4 sch_y=56.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W49 N$98 N$97 "Straight Waveguide" sch_x=-13 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W50 N$100 N$99 "Straight Waveguide" sch_x=-13 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W51 N$102 N$101 "Straight Waveguide" sch_x=-13 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W52 N$104 N$103 "Straight Waveguide" sch_x=-13 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W53 N$106 N$105 "Straight Waveguide" sch_x=-13 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W54 N$108 N$107 "Straight Waveguide" sch_x=-13 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W55 N$110 N$109 "Straight Waveguide" sch_x=-11 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W56 N$112 N$111 "Straight Waveguide" sch_x=-11 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W57 N$114 N$113 "Straight Waveguide" sch_x=-11 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W58 N$116 N$115 "Straight Waveguide" sch_x=-11 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W59 N$118 N$117 "Straight Waveguide" sch_x=-9 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W60 N$120 N$119 "Straight Waveguide" sch_x=-9 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W61 N$121 N$122 "Straight Waveguide" sch_x=-9 sch_y=62.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W62 N$123 N$124 "Straight Waveguide" sch_x=-8 sch_y=61.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W63 N$125 N$126 "Straight Waveguide" sch_x=-7 sch_y=60.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W64 N$127 N$128 "Straight Waveguide" sch_x=-7 sch_y=59.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W65 N$129 N$130 "Straight Waveguide" sch_x=-8 sch_y=58.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W66 N$131 N$132 "Straight Waveguide" sch_x=-9 sch_y=57.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W67 N$133 N$134 "Straight Waveguide" sch_x=-10 sch_y=62.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W68 N$135 N$136 "Straight Waveguide" sch_x=-10 sch_y=57.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W69 N$137 N$138 "Straight Waveguide" sch_x=13 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W70 N$139 N$140 "Straight Waveguide" sch_x=13 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W71 N$141 N$142 "Straight Waveguide" sch_x=13 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W72 N$143 N$144 "Straight Waveguide" sch_x=13 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W73 N$145 N$146 "Straight Waveguide" sch_x=13 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W74 N$147 N$148 "Straight Waveguide" sch_x=13 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W75 N$149 N$150 "Straight Waveguide" sch_x=11 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W76 N$151 N$152 "Straight Waveguide" sch_x=11 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W77 N$153 N$154 "Straight Waveguide" sch_x=11 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W78 N$155 N$156 "Straight Waveguide" sch_x=11 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W79 N$157 N$158 "Straight Waveguide" sch_x=9 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W80 N$159 N$160 "Straight Waveguide" sch_x=9 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W81 N$162 N$161 "Straight Waveguide" sch_x=9 sch_y=62.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W82 N$164 N$163 "Straight Waveguide" sch_x=8 sch_y=61.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W83 N$166 N$165 "Straight Waveguide" sch_x=7 sch_y=60.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W84 N$168 N$167 "Straight Waveguide" sch_x=7 sch_y=59.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W85 N$170 N$169 "Straight Waveguide" sch_x=8 sch_y=58.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W86 N$172 N$171 "Straight Waveguide" sch_x=9 sch_y=57.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W87 N$174 N$173 "Straight Waveguide" sch_x=10 sch_y=62.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W88 N$176 N$175 "Straight Waveguide" sch_x=10 sch_y=57.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W89 N$177 N$178 "Straight Waveguide" sch_x=-4 sch_y=55.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W90 N$179 N$180 "Straight Waveguide" sch_x=-5 sch_y=54.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W91 N$181 N$182 "Straight Waveguide" sch_x=-5 sch_y=53.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W92 N$183 N$184 "Straight Waveguide" sch_x=-3 sch_y=54.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W93 N$185 N$186 "Straight Waveguide" sch_x=-3 sch_y=53.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W94 N$187 N$188 "Straight Waveguide" sch_x=-4 sch_y=52.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W95 N$189 N$190 "Straight Waveguide" sch_x=0 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W96 N$191 N$192 "Straight Waveguide" sch_x=-1 sch_y=55.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W97 N$193 N$194 "Straight Waveguide" sch_x=-1 sch_y=54.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W98 N$195 N$196 "Straight Waveguide" sch_x=1 sch_y=54.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W99 N$197 N$198 "Straight Waveguide" sch_x=1 sch_y=55.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W100 N$199 N$200 "Straight Waveguide" sch_x=0 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W101 N$201 N$202 "Straight Waveguide" sch_x=0 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W102 N$203 N$204 "Straight Waveguide" sch_x=-1 sch_y=53.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W103 N$205 N$206 "Straight Waveguide" sch_x=-1 sch_y=52.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W104 N$207 N$208 "Straight Waveguide" sch_x=1 sch_y=52.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W105 N$209 N$210 "Straight Waveguide" sch_x=1 sch_y=53.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W106 N$211 N$212 "Straight Waveguide" sch_x=0 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W107 N$213 N$214 "Straight Waveguide" sch_x=4 sch_y=55.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W108 N$215 N$216 "Straight Waveguide" sch_x=3 sch_y=54.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W109 N$217 N$218 "Straight Waveguide" sch_x=3 sch_y=53.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W110 N$219 N$220 "Straight Waveguide" sch_x=5 sch_y=53.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W111 N$221 N$222 "Straight Waveguide" sch_x=5 sch_y=54.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W112 N$223 N$224 "Straight Waveguide" sch_x=4 sch_y=52.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W113 N$225 N$226 "Straight Waveguide" sch_x=-4 sch_y=51.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W114 N$227 N$228 "Straight Waveguide" sch_x=-5 sch_y=50.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W115 N$229 N$230 "Straight Waveguide" sch_x=-5 sch_y=49.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W116 N$231 N$232 "Straight Waveguide" sch_x=-3 sch_y=50.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W117 N$233 N$234 "Straight Waveguide" sch_x=-3 sch_y=49.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W118 N$235 N$236 "Straight Waveguide" sch_x=-4 sch_y=48.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W119 N$237 N$238 "Straight Waveguide" sch_x=0 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W120 N$239 N$240 "Straight Waveguide" sch_x=-1 sch_y=51.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W121 N$241 N$242 "Straight Waveguide" sch_x=-1 sch_y=50.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W122 N$243 N$244 "Straight Waveguide" sch_x=1 sch_y=50.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W123 N$245 N$246 "Straight Waveguide" sch_x=1 sch_y=51.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W124 N$247 N$248 "Straight Waveguide" sch_x=0 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W125 N$249 N$250 "Straight Waveguide" sch_x=0 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W126 N$251 N$252 "Straight Waveguide" sch_x=-1 sch_y=49.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W127 N$253 N$254 "Straight Waveguide" sch_x=-1 sch_y=48.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W128 N$255 N$256 "Straight Waveguide" sch_x=1 sch_y=48.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W129 N$257 N$258 "Straight Waveguide" sch_x=1 sch_y=49.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W130 N$259 N$260 "Straight Waveguide" sch_x=0 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W131 N$261 N$262 "Straight Waveguide" sch_x=4 sch_y=51.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W132 N$263 N$264 "Straight Waveguide" sch_x=3 sch_y=50.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W133 N$265 N$266 "Straight Waveguide" sch_x=3 sch_y=49.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W134 N$267 N$268 "Straight Waveguide" sch_x=5 sch_y=49.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W135 N$269 N$270 "Straight Waveguide" sch_x=5 sch_y=50.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W136 N$271 N$272 "Straight Waveguide" sch_x=4 sch_y=48.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W137 N$274 N$273 "Straight Waveguide" sch_x=-13 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W138 N$276 N$275 "Straight Waveguide" sch_x=-13 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W139 N$278 N$277 "Straight Waveguide" sch_x=-13 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W140 N$280 N$279 "Straight Waveguide" sch_x=-13 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W141 N$282 N$281 "Straight Waveguide" sch_x=-13 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W142 N$284 N$283 "Straight Waveguide" sch_x=-13 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W143 N$286 N$285 "Straight Waveguide" sch_x=-11 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W144 N$288 N$287 "Straight Waveguide" sch_x=-11 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W145 N$290 N$289 "Straight Waveguide" sch_x=-11 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W146 N$292 N$291 "Straight Waveguide" sch_x=-11 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W147 N$294 N$293 "Straight Waveguide" sch_x=-9 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W148 N$296 N$295 "Straight Waveguide" sch_x=-9 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W149 N$297 N$298 "Straight Waveguide" sch_x=-9 sch_y=54.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W150 N$299 N$300 "Straight Waveguide" sch_x=-8 sch_y=53.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W151 N$301 N$302 "Straight Waveguide" sch_x=-7 sch_y=52.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W152 N$303 N$304 "Straight Waveguide" sch_x=-7 sch_y=51.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W153 N$305 N$306 "Straight Waveguide" sch_x=-8 sch_y=50.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W154 N$307 N$308 "Straight Waveguide" sch_x=-9 sch_y=49.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W155 N$309 N$310 "Straight Waveguide" sch_x=-10 sch_y=54.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W156 N$311 N$312 "Straight Waveguide" sch_x=-10 sch_y=49.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W157 N$313 N$314 "Straight Waveguide" sch_x=13 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W158 N$315 N$316 "Straight Waveguide" sch_x=13 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W159 N$317 N$318 "Straight Waveguide" sch_x=13 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W160 N$319 N$320 "Straight Waveguide" sch_x=13 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W161 N$321 N$322 "Straight Waveguide" sch_x=13 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W162 N$323 N$324 "Straight Waveguide" sch_x=13 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W163 N$325 N$326 "Straight Waveguide" sch_x=11 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W164 N$327 N$328 "Straight Waveguide" sch_x=11 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W165 N$329 N$330 "Straight Waveguide" sch_x=11 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W166 N$331 N$332 "Straight Waveguide" sch_x=11 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W167 N$333 N$334 "Straight Waveguide" sch_x=9 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W168 N$335 N$336 "Straight Waveguide" sch_x=9 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W169 N$338 N$337 "Straight Waveguide" sch_x=9 sch_y=54.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W170 N$340 N$339 "Straight Waveguide" sch_x=8 sch_y=53.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W171 N$342 N$341 "Straight Waveguide" sch_x=7 sch_y=52.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W172 N$344 N$343 "Straight Waveguide" sch_x=7 sch_y=51.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W173 N$346 N$345 "Straight Waveguide" sch_x=8 sch_y=50.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W174 N$348 N$347 "Straight Waveguide" sch_x=9 sch_y=49.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W175 N$350 N$349 "Straight Waveguide" sch_x=10 sch_y=54.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W176 N$352 N$351 "Straight Waveguide" sch_x=10 sch_y=49.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W177 N$354 N$353 "Straight Waveguide" sch_x=-29 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W178 N$356 N$355 "Straight Waveguide" sch_x=-29 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W179 N$358 N$357 "Straight Waveguide" sch_x=-29 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W180 N$360 N$359 "Straight Waveguide" sch_x=-29 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W181 N$362 N$361 "Straight Waveguide" sch_x=-29 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W182 N$364 N$363 "Straight Waveguide" sch_x=-29 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W183 N$366 N$365 "Straight Waveguide" sch_x=-29 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W184 N$368 N$367 "Straight Waveguide" sch_x=-29 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W185 N$370 N$369 "Straight Waveguide" sch_x=-29 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W186 N$372 N$371 "Straight Waveguide" sch_x=-29 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W187 N$374 N$373 "Straight Waveguide" sch_x=-29 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W188 N$376 N$375 "Straight Waveguide" sch_x=-29 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W189 N$378 N$377 "Straight Waveguide" sch_x=-29 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W190 N$380 N$379 "Straight Waveguide" sch_x=-29 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W191 N$382 N$381 "Straight Waveguide" sch_x=-27 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W192 N$384 N$383 "Straight Waveguide" sch_x=-27 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W193 N$386 N$385 "Straight Waveguide" sch_x=-27 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W194 N$388 N$387 "Straight Waveguide" sch_x=-27 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W195 N$390 N$389 "Straight Waveguide" sch_x=-27 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W196 N$392 N$391 "Straight Waveguide" sch_x=-27 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W197 N$394 N$393 "Straight Waveguide" sch_x=-27 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W198 N$396 N$395 "Straight Waveguide" sch_x=-27 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W199 N$398 N$397 "Straight Waveguide" sch_x=-27 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W200 N$400 N$399 "Straight Waveguide" sch_x=-27 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W201 N$402 N$401 "Straight Waveguide" sch_x=-27 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W202 N$404 N$403 "Straight Waveguide" sch_x=-27 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W203 N$406 N$405 "Straight Waveguide" sch_x=-25 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W204 N$408 N$407 "Straight Waveguide" sch_x=-25 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W205 N$410 N$409 "Straight Waveguide" sch_x=-25 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W206 N$412 N$411 "Straight Waveguide" sch_x=-25 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W207 N$414 N$413 "Straight Waveguide" sch_x=-25 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W208 N$416 N$415 "Straight Waveguide" sch_x=-25 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W209 N$418 N$417 "Straight Waveguide" sch_x=-25 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W210 N$420 N$419 "Straight Waveguide" sch_x=-25 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W211 N$422 N$421 "Straight Waveguide" sch_x=-25 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W212 N$424 N$423 "Straight Waveguide" sch_x=-25 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W213 N$426 N$425 "Straight Waveguide" sch_x=-23 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W214 N$428 N$427 "Straight Waveguide" sch_x=-23 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W215 N$430 N$429 "Straight Waveguide" sch_x=-23 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W216 N$432 N$431 "Straight Waveguide" sch_x=-23 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W217 N$434 N$433 "Straight Waveguide" sch_x=-23 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W218 N$436 N$435 "Straight Waveguide" sch_x=-23 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W219 N$438 N$437 "Straight Waveguide" sch_x=-23 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W220 N$440 N$439 "Straight Waveguide" sch_x=-23 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W221 N$442 N$441 "Straight Waveguide" sch_x=-21 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W222 N$444 N$443 "Straight Waveguide" sch_x=-21 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W223 N$446 N$445 "Straight Waveguide" sch_x=-21 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W224 N$448 N$447 "Straight Waveguide" sch_x=-21 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W225 N$450 N$449 "Straight Waveguide" sch_x=-21 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W226 N$452 N$451 "Straight Waveguide" sch_x=-21 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W227 N$454 N$453 "Straight Waveguide" sch_x=-19 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W228 N$456 N$455 "Straight Waveguide" sch_x=-19 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W229 N$458 N$457 "Straight Waveguide" sch_x=-19 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W230 N$460 N$459 "Straight Waveguide" sch_x=-19 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W231 N$462 N$461 "Straight Waveguide" sch_x=-17 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W232 N$464 N$463 "Straight Waveguide" sch_x=-17 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W233 N$465 N$466 "Straight Waveguide" sch_x=-21 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W234 N$467 N$468 "Straight Waveguide" sch_x=-20 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W235 N$469 N$470 "Straight Waveguide" sch_x=-19 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W236 N$471 N$472 "Straight Waveguide" sch_x=-18 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W237 N$473 N$474 "Straight Waveguide" sch_x=-17 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W238 N$475 N$476 "Straight Waveguide" sch_x=-16 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W239 N$477 N$478 "Straight Waveguide" sch_x=-15 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W240 N$479 N$480 "Straight Waveguide" sch_x=-15 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W241 N$481 N$482 "Straight Waveguide" sch_x=-16 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W242 N$483 N$484 "Straight Waveguide" sch_x=-17 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W243 N$485 N$486 "Straight Waveguide" sch_x=-18 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W244 N$487 N$488 "Straight Waveguide" sch_x=-19 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W245 N$489 N$490 "Straight Waveguide" sch_x=-20 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W246 N$491 N$492 "Straight Waveguide" sch_x=-21 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W247 N$493 N$494 "Straight Waveguide" sch_x=-22 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W248 N$495 N$496 "Straight Waveguide" sch_x=-22 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W249 N$497 N$498 "Straight Waveguide" sch_x=29 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W250 N$499 N$500 "Straight Waveguide" sch_x=29 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W251 N$501 N$502 "Straight Waveguide" sch_x=29 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W252 N$503 N$504 "Straight Waveguide" sch_x=29 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W253 N$505 N$506 "Straight Waveguide" sch_x=29 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W254 N$507 N$508 "Straight Waveguide" sch_x=29 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W255 N$509 N$510 "Straight Waveguide" sch_x=29 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W256 N$511 N$512 "Straight Waveguide" sch_x=29 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W257 N$513 N$514 "Straight Waveguide" sch_x=29 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W258 N$515 N$516 "Straight Waveguide" sch_x=29 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W259 N$517 N$518 "Straight Waveguide" sch_x=29 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W260 N$519 N$520 "Straight Waveguide" sch_x=29 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W261 N$521 N$522 "Straight Waveguide" sch_x=29 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W262 N$523 N$524 "Straight Waveguide" sch_x=29 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W263 N$525 N$526 "Straight Waveguide" sch_x=27 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W264 N$527 N$528 "Straight Waveguide" sch_x=27 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W265 N$529 N$530 "Straight Waveguide" sch_x=27 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W266 N$531 N$532 "Straight Waveguide" sch_x=27 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W267 N$533 N$534 "Straight Waveguide" sch_x=27 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W268 N$535 N$536 "Straight Waveguide" sch_x=27 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W269 N$537 N$538 "Straight Waveguide" sch_x=27 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W270 N$539 N$540 "Straight Waveguide" sch_x=27 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W271 N$541 N$542 "Straight Waveguide" sch_x=27 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W272 N$543 N$544 "Straight Waveguide" sch_x=27 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W273 N$545 N$546 "Straight Waveguide" sch_x=27 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W274 N$547 N$548 "Straight Waveguide" sch_x=27 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W275 N$549 N$550 "Straight Waveguide" sch_x=25 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W276 N$551 N$552 "Straight Waveguide" sch_x=25 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W277 N$553 N$554 "Straight Waveguide" sch_x=25 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W278 N$555 N$556 "Straight Waveguide" sch_x=25 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W279 N$557 N$558 "Straight Waveguide" sch_x=25 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W280 N$559 N$560 "Straight Waveguide" sch_x=25 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W281 N$561 N$562 "Straight Waveguide" sch_x=25 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W282 N$563 N$564 "Straight Waveguide" sch_x=25 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W283 N$565 N$566 "Straight Waveguide" sch_x=25 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W284 N$567 N$568 "Straight Waveguide" sch_x=25 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W285 N$569 N$570 "Straight Waveguide" sch_x=23 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W286 N$571 N$572 "Straight Waveguide" sch_x=23 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W287 N$573 N$574 "Straight Waveguide" sch_x=23 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W288 N$575 N$576 "Straight Waveguide" sch_x=23 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W289 N$577 N$578 "Straight Waveguide" sch_x=23 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W290 N$579 N$580 "Straight Waveguide" sch_x=23 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W291 N$581 N$582 "Straight Waveguide" sch_x=23 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W292 N$583 N$584 "Straight Waveguide" sch_x=23 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W293 N$585 N$586 "Straight Waveguide" sch_x=21 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W294 N$587 N$588 "Straight Waveguide" sch_x=21 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W295 N$589 N$590 "Straight Waveguide" sch_x=21 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W296 N$591 N$592 "Straight Waveguide" sch_x=21 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W297 N$593 N$594 "Straight Waveguide" sch_x=21 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W298 N$595 N$596 "Straight Waveguide" sch_x=21 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W299 N$597 N$598 "Straight Waveguide" sch_x=19 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W300 N$599 N$600 "Straight Waveguide" sch_x=19 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W301 N$601 N$602 "Straight Waveguide" sch_x=19 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W302 N$603 N$604 "Straight Waveguide" sch_x=19 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W303 N$605 N$606 "Straight Waveguide" sch_x=17 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W304 N$607 N$608 "Straight Waveguide" sch_x=17 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W305 N$610 N$609 "Straight Waveguide" sch_x=21 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W306 N$612 N$611 "Straight Waveguide" sch_x=20 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W307 N$614 N$613 "Straight Waveguide" sch_x=19 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W308 N$616 N$615 "Straight Waveguide" sch_x=18 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W309 N$618 N$617 "Straight Waveguide" sch_x=17 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W310 N$620 N$619 "Straight Waveguide" sch_x=16 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W311 N$622 N$621 "Straight Waveguide" sch_x=15 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W312 N$624 N$623 "Straight Waveguide" sch_x=15 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W313 N$626 N$625 "Straight Waveguide" sch_x=16 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W314 N$628 N$627 "Straight Waveguide" sch_x=17 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W315 N$630 N$629 "Straight Waveguide" sch_x=18 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W316 N$632 N$631 "Straight Waveguide" sch_x=19 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W317 N$634 N$633 "Straight Waveguide" sch_x=20 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W318 N$636 N$635 "Straight Waveguide" sch_x=21 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W319 N$638 N$637 "Straight Waveguide" sch_x=22 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W320 N$640 N$639 "Straight Waveguide" sch_x=22 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W321 N$641 N$642 "Straight Waveguide" sch_x=-4 sch_y=47.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W322 N$643 N$644 "Straight Waveguide" sch_x=-5 sch_y=46.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W323 N$645 N$646 "Straight Waveguide" sch_x=-5 sch_y=45.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W324 N$647 N$648 "Straight Waveguide" sch_x=-3 sch_y=46.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W325 N$649 N$650 "Straight Waveguide" sch_x=-3 sch_y=45.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W326 N$651 N$652 "Straight Waveguide" sch_x=-4 sch_y=44.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W327 N$653 N$654 "Straight Waveguide" sch_x=0 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W328 N$655 N$656 "Straight Waveguide" sch_x=-1 sch_y=47.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W329 N$657 N$658 "Straight Waveguide" sch_x=-1 sch_y=46.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W330 N$659 N$660 "Straight Waveguide" sch_x=1 sch_y=46.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W331 N$661 N$662 "Straight Waveguide" sch_x=1 sch_y=47.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W332 N$663 N$664 "Straight Waveguide" sch_x=0 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W333 N$665 N$666 "Straight Waveguide" sch_x=0 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W334 N$667 N$668 "Straight Waveguide" sch_x=-1 sch_y=45.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W335 N$669 N$670 "Straight Waveguide" sch_x=-1 sch_y=44.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W336 N$671 N$672 "Straight Waveguide" sch_x=1 sch_y=44.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W337 N$673 N$674 "Straight Waveguide" sch_x=1 sch_y=45.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W338 N$675 N$676 "Straight Waveguide" sch_x=0 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W339 N$677 N$678 "Straight Waveguide" sch_x=4 sch_y=47.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W340 N$679 N$680 "Straight Waveguide" sch_x=3 sch_y=46.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W341 N$681 N$682 "Straight Waveguide" sch_x=3 sch_y=45.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W342 N$683 N$684 "Straight Waveguide" sch_x=5 sch_y=45.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W343 N$685 N$686 "Straight Waveguide" sch_x=5 sch_y=46.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W344 N$687 N$688 "Straight Waveguide" sch_x=4 sch_y=44.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W345 N$689 N$690 "Straight Waveguide" sch_x=-4 sch_y=43.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W346 N$691 N$692 "Straight Waveguide" sch_x=-5 sch_y=42.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W347 N$693 N$694 "Straight Waveguide" sch_x=-5 sch_y=41.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W348 N$695 N$696 "Straight Waveguide" sch_x=-3 sch_y=42.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W349 N$697 N$698 "Straight Waveguide" sch_x=-3 sch_y=41.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W350 N$699 N$700 "Straight Waveguide" sch_x=-4 sch_y=40.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W351 N$701 N$702 "Straight Waveguide" sch_x=0 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W352 N$703 N$704 "Straight Waveguide" sch_x=-1 sch_y=43.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W353 N$705 N$706 "Straight Waveguide" sch_x=-1 sch_y=42.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W354 N$707 N$708 "Straight Waveguide" sch_x=1 sch_y=42.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W355 N$709 N$710 "Straight Waveguide" sch_x=1 sch_y=43.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W356 N$711 N$712 "Straight Waveguide" sch_x=0 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W357 N$713 N$714 "Straight Waveguide" sch_x=0 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W358 N$715 N$716 "Straight Waveguide" sch_x=-1 sch_y=41.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W359 N$717 N$718 "Straight Waveguide" sch_x=-1 sch_y=40.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W360 N$719 N$720 "Straight Waveguide" sch_x=1 sch_y=40.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W361 N$721 N$722 "Straight Waveguide" sch_x=1 sch_y=41.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W362 N$723 N$724 "Straight Waveguide" sch_x=0 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W363 N$725 N$726 "Straight Waveguide" sch_x=4 sch_y=43.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W364 N$727 N$728 "Straight Waveguide" sch_x=3 sch_y=42.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W365 N$729 N$730 "Straight Waveguide" sch_x=3 sch_y=41.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W366 N$731 N$732 "Straight Waveguide" sch_x=5 sch_y=41.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W367 N$733 N$734 "Straight Waveguide" sch_x=5 sch_y=42.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W368 N$735 N$736 "Straight Waveguide" sch_x=4 sch_y=40.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W369 N$738 N$737 "Straight Waveguide" sch_x=-13 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W370 N$740 N$739 "Straight Waveguide" sch_x=-13 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W371 N$742 N$741 "Straight Waveguide" sch_x=-13 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W372 N$744 N$743 "Straight Waveguide" sch_x=-13 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W373 N$746 N$745 "Straight Waveguide" sch_x=-13 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W374 N$748 N$747 "Straight Waveguide" sch_x=-13 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W375 N$750 N$749 "Straight Waveguide" sch_x=-11 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W376 N$752 N$751 "Straight Waveguide" sch_x=-11 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W377 N$754 N$753 "Straight Waveguide" sch_x=-11 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W378 N$756 N$755 "Straight Waveguide" sch_x=-11 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W379 N$758 N$757 "Straight Waveguide" sch_x=-9 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W380 N$760 N$759 "Straight Waveguide" sch_x=-9 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W381 N$761 N$762 "Straight Waveguide" sch_x=-9 sch_y=46.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W382 N$763 N$764 "Straight Waveguide" sch_x=-8 sch_y=45.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W383 N$765 N$766 "Straight Waveguide" sch_x=-7 sch_y=44.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W384 N$767 N$768 "Straight Waveguide" sch_x=-7 sch_y=43.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W385 N$769 N$770 "Straight Waveguide" sch_x=-8 sch_y=42.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W386 N$771 N$772 "Straight Waveguide" sch_x=-9 sch_y=41.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W387 N$773 N$774 "Straight Waveguide" sch_x=-10 sch_y=46.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W388 N$775 N$776 "Straight Waveguide" sch_x=-10 sch_y=41.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W389 N$777 N$778 "Straight Waveguide" sch_x=13 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W390 N$779 N$780 "Straight Waveguide" sch_x=13 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W391 N$781 N$782 "Straight Waveguide" sch_x=13 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W392 N$783 N$784 "Straight Waveguide" sch_x=13 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W393 N$785 N$786 "Straight Waveguide" sch_x=13 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W394 N$787 N$788 "Straight Waveguide" sch_x=13 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W395 N$789 N$790 "Straight Waveguide" sch_x=11 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W396 N$791 N$792 "Straight Waveguide" sch_x=11 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W397 N$793 N$794 "Straight Waveguide" sch_x=11 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W398 N$795 N$796 "Straight Waveguide" sch_x=11 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W399 N$797 N$798 "Straight Waveguide" sch_x=9 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W400 N$799 N$800 "Straight Waveguide" sch_x=9 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W401 N$802 N$801 "Straight Waveguide" sch_x=9 sch_y=46.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W402 N$804 N$803 "Straight Waveguide" sch_x=8 sch_y=45.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W403 N$806 N$805 "Straight Waveguide" sch_x=7 sch_y=44.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W404 N$808 N$807 "Straight Waveguide" sch_x=7 sch_y=43.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W405 N$810 N$809 "Straight Waveguide" sch_x=8 sch_y=42.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W406 N$812 N$811 "Straight Waveguide" sch_x=9 sch_y=41.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W407 N$814 N$813 "Straight Waveguide" sch_x=10 sch_y=46.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W408 N$816 N$815 "Straight Waveguide" sch_x=10 sch_y=41.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W409 N$817 N$818 "Straight Waveguide" sch_x=-4 sch_y=39.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W410 N$819 N$820 "Straight Waveguide" sch_x=-5 sch_y=38.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W411 N$821 N$822 "Straight Waveguide" sch_x=-5 sch_y=37.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W412 N$823 N$824 "Straight Waveguide" sch_x=-3 sch_y=38.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W413 N$825 N$826 "Straight Waveguide" sch_x=-3 sch_y=37.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W414 N$827 N$828 "Straight Waveguide" sch_x=-4 sch_y=36.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W415 N$829 N$830 "Straight Waveguide" sch_x=0 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W416 N$831 N$832 "Straight Waveguide" sch_x=-1 sch_y=39.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W417 N$833 N$834 "Straight Waveguide" sch_x=-1 sch_y=38.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W418 N$835 N$836 "Straight Waveguide" sch_x=1 sch_y=38.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W419 N$837 N$838 "Straight Waveguide" sch_x=1 sch_y=39.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W420 N$839 N$840 "Straight Waveguide" sch_x=0 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W421 N$841 N$842 "Straight Waveguide" sch_x=0 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W422 N$843 N$844 "Straight Waveguide" sch_x=-1 sch_y=37.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W423 N$845 N$846 "Straight Waveguide" sch_x=-1 sch_y=36.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W424 N$847 N$848 "Straight Waveguide" sch_x=1 sch_y=36.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W425 N$849 N$850 "Straight Waveguide" sch_x=1 sch_y=37.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W426 N$851 N$852 "Straight Waveguide" sch_x=0 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W427 N$853 N$854 "Straight Waveguide" sch_x=4 sch_y=39.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W428 N$855 N$856 "Straight Waveguide" sch_x=3 sch_y=38.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W429 N$857 N$858 "Straight Waveguide" sch_x=3 sch_y=37.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W430 N$859 N$860 "Straight Waveguide" sch_x=5 sch_y=37.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W431 N$861 N$862 "Straight Waveguide" sch_x=5 sch_y=38.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W432 N$863 N$864 "Straight Waveguide" sch_x=4 sch_y=36.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W433 N$865 N$866 "Straight Waveguide" sch_x=-4 sch_y=35.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W434 N$867 N$868 "Straight Waveguide" sch_x=-5 sch_y=34.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W435 N$869 N$870 "Straight Waveguide" sch_x=-5 sch_y=33.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W436 N$871 N$872 "Straight Waveguide" sch_x=-3 sch_y=34.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W437 N$873 N$874 "Straight Waveguide" sch_x=-3 sch_y=33.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W438 N$875 N$876 "Straight Waveguide" sch_x=-4 sch_y=32.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W439 N$877 N$878 "Straight Waveguide" sch_x=0 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W440 N$879 N$880 "Straight Waveguide" sch_x=-1 sch_y=35.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W441 N$881 N$882 "Straight Waveguide" sch_x=-1 sch_y=34.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W442 N$883 N$884 "Straight Waveguide" sch_x=1 sch_y=34.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W443 N$885 N$886 "Straight Waveguide" sch_x=1 sch_y=35.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W444 N$887 N$888 "Straight Waveguide" sch_x=0 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W445 N$889 N$890 "Straight Waveguide" sch_x=0 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W446 N$891 N$892 "Straight Waveguide" sch_x=-1 sch_y=33.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W447 N$893 N$894 "Straight Waveguide" sch_x=-1 sch_y=32.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W448 N$895 N$896 "Straight Waveguide" sch_x=1 sch_y=32.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W449 N$897 N$898 "Straight Waveguide" sch_x=1 sch_y=33.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W450 N$899 N$900 "Straight Waveguide" sch_x=0 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W451 N$901 N$902 "Straight Waveguide" sch_x=4 sch_y=35.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W452 N$903 N$904 "Straight Waveguide" sch_x=3 sch_y=34.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W453 N$905 N$906 "Straight Waveguide" sch_x=3 sch_y=33.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W454 N$907 N$908 "Straight Waveguide" sch_x=5 sch_y=33.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W455 N$909 N$910 "Straight Waveguide" sch_x=5 sch_y=34.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W456 N$911 N$912 "Straight Waveguide" sch_x=4 sch_y=32.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W457 N$914 N$913 "Straight Waveguide" sch_x=-13 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W458 N$916 N$915 "Straight Waveguide" sch_x=-13 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W459 N$918 N$917 "Straight Waveguide" sch_x=-13 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W460 N$920 N$919 "Straight Waveguide" sch_x=-13 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W461 N$922 N$921 "Straight Waveguide" sch_x=-13 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W462 N$924 N$923 "Straight Waveguide" sch_x=-13 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W463 N$926 N$925 "Straight Waveguide" sch_x=-11 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W464 N$928 N$927 "Straight Waveguide" sch_x=-11 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W465 N$930 N$929 "Straight Waveguide" sch_x=-11 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W466 N$932 N$931 "Straight Waveguide" sch_x=-11 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W467 N$934 N$933 "Straight Waveguide" sch_x=-9 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W468 N$936 N$935 "Straight Waveguide" sch_x=-9 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W469 N$937 N$938 "Straight Waveguide" sch_x=-9 sch_y=38.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W470 N$939 N$940 "Straight Waveguide" sch_x=-8 sch_y=37.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W471 N$941 N$942 "Straight Waveguide" sch_x=-7 sch_y=36.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W472 N$943 N$944 "Straight Waveguide" sch_x=-7 sch_y=35.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W473 N$945 N$946 "Straight Waveguide" sch_x=-8 sch_y=34.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W474 N$947 N$948 "Straight Waveguide" sch_x=-9 sch_y=33.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W475 N$949 N$950 "Straight Waveguide" sch_x=-10 sch_y=38.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W476 N$951 N$952 "Straight Waveguide" sch_x=-10 sch_y=33.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W477 N$953 N$954 "Straight Waveguide" sch_x=13 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W478 N$955 N$956 "Straight Waveguide" sch_x=13 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W479 N$957 N$958 "Straight Waveguide" sch_x=13 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W480 N$959 N$960 "Straight Waveguide" sch_x=13 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W481 N$961 N$962 "Straight Waveguide" sch_x=13 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W482 N$963 N$964 "Straight Waveguide" sch_x=13 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W483 N$965 N$966 "Straight Waveguide" sch_x=11 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W484 N$967 N$968 "Straight Waveguide" sch_x=11 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W485 N$969 N$970 "Straight Waveguide" sch_x=11 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W486 N$971 N$972 "Straight Waveguide" sch_x=11 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W487 N$973 N$974 "Straight Waveguide" sch_x=9 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W488 N$975 N$976 "Straight Waveguide" sch_x=9 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W489 N$978 N$977 "Straight Waveguide" sch_x=9 sch_y=38.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W490 N$980 N$979 "Straight Waveguide" sch_x=8 sch_y=37.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W491 N$982 N$981 "Straight Waveguide" sch_x=7 sch_y=36.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W492 N$984 N$983 "Straight Waveguide" sch_x=7 sch_y=35.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W493 N$986 N$985 "Straight Waveguide" sch_x=8 sch_y=34.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W494 N$988 N$987 "Straight Waveguide" sch_x=9 sch_y=33.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W495 N$990 N$989 "Straight Waveguide" sch_x=10 sch_y=38.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W496 N$992 N$991 "Straight Waveguide" sch_x=10 sch_y=33.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W497 N$994 N$993 "Straight Waveguide" sch_x=-29 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W498 N$996 N$995 "Straight Waveguide" sch_x=-29 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W499 N$998 N$997 "Straight Waveguide" sch_x=-29 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W500 N$1000 N$999 "Straight Waveguide" sch_x=-29 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W501 N$1002 N$1001 "Straight Waveguide" sch_x=-29 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W502 N$1004 N$1003 "Straight Waveguide" sch_x=-29 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W503 N$1006 N$1005 "Straight Waveguide" sch_x=-29 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W504 N$1008 N$1007 "Straight Waveguide" sch_x=-29 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W505 N$1010 N$1009 "Straight Waveguide" sch_x=-29 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W506 N$1012 N$1011 "Straight Waveguide" sch_x=-29 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W507 N$1014 N$1013 "Straight Waveguide" sch_x=-29 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W508 N$1016 N$1015 "Straight Waveguide" sch_x=-29 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W509 N$1018 N$1017 "Straight Waveguide" sch_x=-29 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W510 N$1020 N$1019 "Straight Waveguide" sch_x=-29 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W511 N$1022 N$1021 "Straight Waveguide" sch_x=-27 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W512 N$1024 N$1023 "Straight Waveguide" sch_x=-27 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W513 N$1026 N$1025 "Straight Waveguide" sch_x=-27 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W514 N$1028 N$1027 "Straight Waveguide" sch_x=-27 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W515 N$1030 N$1029 "Straight Waveguide" sch_x=-27 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W516 N$1032 N$1031 "Straight Waveguide" sch_x=-27 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W517 N$1034 N$1033 "Straight Waveguide" sch_x=-27 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W518 N$1036 N$1035 "Straight Waveguide" sch_x=-27 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W519 N$1038 N$1037 "Straight Waveguide" sch_x=-27 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W520 N$1040 N$1039 "Straight Waveguide" sch_x=-27 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W521 N$1042 N$1041 "Straight Waveguide" sch_x=-27 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W522 N$1044 N$1043 "Straight Waveguide" sch_x=-27 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W523 N$1046 N$1045 "Straight Waveguide" sch_x=-25 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W524 N$1048 N$1047 "Straight Waveguide" sch_x=-25 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W525 N$1050 N$1049 "Straight Waveguide" sch_x=-25 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W526 N$1052 N$1051 "Straight Waveguide" sch_x=-25 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W527 N$1054 N$1053 "Straight Waveguide" sch_x=-25 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W528 N$1056 N$1055 "Straight Waveguide" sch_x=-25 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W529 N$1058 N$1057 "Straight Waveguide" sch_x=-25 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W530 N$1060 N$1059 "Straight Waveguide" sch_x=-25 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W531 N$1062 N$1061 "Straight Waveguide" sch_x=-25 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W532 N$1064 N$1063 "Straight Waveguide" sch_x=-25 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W533 N$1066 N$1065 "Straight Waveguide" sch_x=-23 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W534 N$1068 N$1067 "Straight Waveguide" sch_x=-23 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W535 N$1070 N$1069 "Straight Waveguide" sch_x=-23 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W536 N$1072 N$1071 "Straight Waveguide" sch_x=-23 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W537 N$1074 N$1073 "Straight Waveguide" sch_x=-23 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W538 N$1076 N$1075 "Straight Waveguide" sch_x=-23 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W539 N$1078 N$1077 "Straight Waveguide" sch_x=-23 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W540 N$1080 N$1079 "Straight Waveguide" sch_x=-23 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W541 N$1082 N$1081 "Straight Waveguide" sch_x=-21 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W542 N$1084 N$1083 "Straight Waveguide" sch_x=-21 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W543 N$1086 N$1085 "Straight Waveguide" sch_x=-21 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W544 N$1088 N$1087 "Straight Waveguide" sch_x=-21 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W545 N$1090 N$1089 "Straight Waveguide" sch_x=-21 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W546 N$1092 N$1091 "Straight Waveguide" sch_x=-21 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W547 N$1094 N$1093 "Straight Waveguide" sch_x=-19 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W548 N$1096 N$1095 "Straight Waveguide" sch_x=-19 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W549 N$1098 N$1097 "Straight Waveguide" sch_x=-19 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W550 N$1100 N$1099 "Straight Waveguide" sch_x=-19 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W551 N$1102 N$1101 "Straight Waveguide" sch_x=-17 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W552 N$1104 N$1103 "Straight Waveguide" sch_x=-17 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W553 N$1105 N$1106 "Straight Waveguide" sch_x=-21 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W554 N$1107 N$1108 "Straight Waveguide" sch_x=-20 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W555 N$1109 N$1110 "Straight Waveguide" sch_x=-19 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W556 N$1111 N$1112 "Straight Waveguide" sch_x=-18 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W557 N$1113 N$1114 "Straight Waveguide" sch_x=-17 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W558 N$1115 N$1116 "Straight Waveguide" sch_x=-16 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W559 N$1117 N$1118 "Straight Waveguide" sch_x=-15 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W560 N$1119 N$1120 "Straight Waveguide" sch_x=-15 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W561 N$1121 N$1122 "Straight Waveguide" sch_x=-16 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W562 N$1123 N$1124 "Straight Waveguide" sch_x=-17 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W563 N$1125 N$1126 "Straight Waveguide" sch_x=-18 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W564 N$1127 N$1128 "Straight Waveguide" sch_x=-19 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W565 N$1129 N$1130 "Straight Waveguide" sch_x=-20 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W566 N$1131 N$1132 "Straight Waveguide" sch_x=-21 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W567 N$1133 N$1134 "Straight Waveguide" sch_x=-22 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W568 N$1135 N$1136 "Straight Waveguide" sch_x=-22 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W569 N$1137 N$1138 "Straight Waveguide" sch_x=29 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W570 N$1139 N$1140 "Straight Waveguide" sch_x=29 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W571 N$1141 N$1142 "Straight Waveguide" sch_x=29 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W572 N$1143 N$1144 "Straight Waveguide" sch_x=29 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W573 N$1145 N$1146 "Straight Waveguide" sch_x=29 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W574 N$1147 N$1148 "Straight Waveguide" sch_x=29 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W575 N$1149 N$1150 "Straight Waveguide" sch_x=29 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W576 N$1151 N$1152 "Straight Waveguide" sch_x=29 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W577 N$1153 N$1154 "Straight Waveguide" sch_x=29 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W578 N$1155 N$1156 "Straight Waveguide" sch_x=29 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W579 N$1157 N$1158 "Straight Waveguide" sch_x=29 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W580 N$1159 N$1160 "Straight Waveguide" sch_x=29 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W581 N$1161 N$1162 "Straight Waveguide" sch_x=29 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W582 N$1163 N$1164 "Straight Waveguide" sch_x=29 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W583 N$1165 N$1166 "Straight Waveguide" sch_x=27 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W584 N$1167 N$1168 "Straight Waveguide" sch_x=27 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W585 N$1169 N$1170 "Straight Waveguide" sch_x=27 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W586 N$1171 N$1172 "Straight Waveguide" sch_x=27 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W587 N$1173 N$1174 "Straight Waveguide" sch_x=27 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W588 N$1175 N$1176 "Straight Waveguide" sch_x=27 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W589 N$1177 N$1178 "Straight Waveguide" sch_x=27 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W590 N$1179 N$1180 "Straight Waveguide" sch_x=27 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W591 N$1181 N$1182 "Straight Waveguide" sch_x=27 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W592 N$1183 N$1184 "Straight Waveguide" sch_x=27 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W593 N$1185 N$1186 "Straight Waveguide" sch_x=27 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W594 N$1187 N$1188 "Straight Waveguide" sch_x=27 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W595 N$1189 N$1190 "Straight Waveguide" sch_x=25 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W596 N$1191 N$1192 "Straight Waveguide" sch_x=25 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W597 N$1193 N$1194 "Straight Waveguide" sch_x=25 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W598 N$1195 N$1196 "Straight Waveguide" sch_x=25 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W599 N$1197 N$1198 "Straight Waveguide" sch_x=25 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W600 N$1199 N$1200 "Straight Waveguide" sch_x=25 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W601 N$1201 N$1202 "Straight Waveguide" sch_x=25 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W602 N$1203 N$1204 "Straight Waveguide" sch_x=25 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W603 N$1205 N$1206 "Straight Waveguide" sch_x=25 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W604 N$1207 N$1208 "Straight Waveguide" sch_x=25 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W605 N$1209 N$1210 "Straight Waveguide" sch_x=23 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W606 N$1211 N$1212 "Straight Waveguide" sch_x=23 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W607 N$1213 N$1214 "Straight Waveguide" sch_x=23 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W608 N$1215 N$1216 "Straight Waveguide" sch_x=23 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W609 N$1217 N$1218 "Straight Waveguide" sch_x=23 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W610 N$1219 N$1220 "Straight Waveguide" sch_x=23 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W611 N$1221 N$1222 "Straight Waveguide" sch_x=23 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W612 N$1223 N$1224 "Straight Waveguide" sch_x=23 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W613 N$1225 N$1226 "Straight Waveguide" sch_x=21 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W614 N$1227 N$1228 "Straight Waveguide" sch_x=21 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W615 N$1229 N$1230 "Straight Waveguide" sch_x=21 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W616 N$1231 N$1232 "Straight Waveguide" sch_x=21 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W617 N$1233 N$1234 "Straight Waveguide" sch_x=21 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W618 N$1235 N$1236 "Straight Waveguide" sch_x=21 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W619 N$1237 N$1238 "Straight Waveguide" sch_x=19 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W620 N$1239 N$1240 "Straight Waveguide" sch_x=19 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W621 N$1241 N$1242 "Straight Waveguide" sch_x=19 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W622 N$1243 N$1244 "Straight Waveguide" sch_x=19 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W623 N$1245 N$1246 "Straight Waveguide" sch_x=17 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W624 N$1247 N$1248 "Straight Waveguide" sch_x=17 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W625 N$1250 N$1249 "Straight Waveguide" sch_x=21 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W626 N$1252 N$1251 "Straight Waveguide" sch_x=20 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W627 N$1254 N$1253 "Straight Waveguide" sch_x=19 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W628 N$1256 N$1255 "Straight Waveguide" sch_x=18 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W629 N$1258 N$1257 "Straight Waveguide" sch_x=17 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W630 N$1260 N$1259 "Straight Waveguide" sch_x=16 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W631 N$1262 N$1261 "Straight Waveguide" sch_x=15 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W632 N$1264 N$1263 "Straight Waveguide" sch_x=15 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W633 N$1266 N$1265 "Straight Waveguide" sch_x=16 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W634 N$1268 N$1267 "Straight Waveguide" sch_x=17 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W635 N$1270 N$1269 "Straight Waveguide" sch_x=18 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W636 N$1272 N$1271 "Straight Waveguide" sch_x=19 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W637 N$1274 N$1273 "Straight Waveguide" sch_x=20 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W638 N$1276 N$1275 "Straight Waveguide" sch_x=21 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W639 N$1278 N$1277 "Straight Waveguide" sch_x=22 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W640 N$1280 N$1279 "Straight Waveguide" sch_x=22 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W641 N$1282 N$1281 "Straight Waveguide" sch_x=-61 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W642 N$1284 N$1283 "Straight Waveguide" sch_x=-61 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W643 N$1286 N$1285 "Straight Waveguide" sch_x=-61 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W644 N$1288 N$1287 "Straight Waveguide" sch_x=-61 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W645 N$1290 N$1289 "Straight Waveguide" sch_x=-61 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W646 N$1292 N$1291 "Straight Waveguide" sch_x=-61 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W647 N$1294 N$1293 "Straight Waveguide" sch_x=-61 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W648 N$1296 N$1295 "Straight Waveguide" sch_x=-61 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W649 N$1298 N$1297 "Straight Waveguide" sch_x=-61 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W650 N$1300 N$1299 "Straight Waveguide" sch_x=-61 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W651 N$1302 N$1301 "Straight Waveguide" sch_x=-61 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W652 N$1304 N$1303 "Straight Waveguide" sch_x=-61 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W653 N$1306 N$1305 "Straight Waveguide" sch_x=-61 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W654 N$1308 N$1307 "Straight Waveguide" sch_x=-61 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W655 N$1310 N$1309 "Straight Waveguide" sch_x=-61 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W656 N$1312 N$1311 "Straight Waveguide" sch_x=-61 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W657 N$1314 N$1313 "Straight Waveguide" sch_x=-61 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W658 N$1316 N$1315 "Straight Waveguide" sch_x=-61 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W659 N$1318 N$1317 "Straight Waveguide" sch_x=-61 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W660 N$1320 N$1319 "Straight Waveguide" sch_x=-61 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W661 N$1322 N$1321 "Straight Waveguide" sch_x=-61 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W662 N$1324 N$1323 "Straight Waveguide" sch_x=-61 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W663 N$1326 N$1325 "Straight Waveguide" sch_x=-61 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W664 N$1328 N$1327 "Straight Waveguide" sch_x=-61 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W665 N$1330 N$1329 "Straight Waveguide" sch_x=-61 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W666 N$1332 N$1331 "Straight Waveguide" sch_x=-61 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W667 N$1334 N$1333 "Straight Waveguide" sch_x=-61 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W668 N$1336 N$1335 "Straight Waveguide" sch_x=-61 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W669 N$1338 N$1337 "Straight Waveguide" sch_x=-61 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W670 N$1340 N$1339 "Straight Waveguide" sch_x=-61 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W671 N$1342 N$1341 "Straight Waveguide" sch_x=-59 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W672 N$1344 N$1343 "Straight Waveguide" sch_x=-59 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W673 N$1346 N$1345 "Straight Waveguide" sch_x=-59 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W674 N$1348 N$1347 "Straight Waveguide" sch_x=-59 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W675 N$1350 N$1349 "Straight Waveguide" sch_x=-59 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W676 N$1352 N$1351 "Straight Waveguide" sch_x=-59 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W677 N$1354 N$1353 "Straight Waveguide" sch_x=-59 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W678 N$1356 N$1355 "Straight Waveguide" sch_x=-59 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W679 N$1358 N$1357 "Straight Waveguide" sch_x=-59 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W680 N$1360 N$1359 "Straight Waveguide" sch_x=-59 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W681 N$1362 N$1361 "Straight Waveguide" sch_x=-59 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W682 N$1364 N$1363 "Straight Waveguide" sch_x=-59 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W683 N$1366 N$1365 "Straight Waveguide" sch_x=-59 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W684 N$1368 N$1367 "Straight Waveguide" sch_x=-59 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W685 N$1370 N$1369 "Straight Waveguide" sch_x=-59 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W686 N$1372 N$1371 "Straight Waveguide" sch_x=-59 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W687 N$1374 N$1373 "Straight Waveguide" sch_x=-59 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W688 N$1376 N$1375 "Straight Waveguide" sch_x=-59 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W689 N$1378 N$1377 "Straight Waveguide" sch_x=-59 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W690 N$1380 N$1379 "Straight Waveguide" sch_x=-59 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W691 N$1382 N$1381 "Straight Waveguide" sch_x=-59 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W692 N$1384 N$1383 "Straight Waveguide" sch_x=-59 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W693 N$1386 N$1385 "Straight Waveguide" sch_x=-59 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W694 N$1388 N$1387 "Straight Waveguide" sch_x=-59 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W695 N$1390 N$1389 "Straight Waveguide" sch_x=-59 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W696 N$1392 N$1391 "Straight Waveguide" sch_x=-59 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W697 N$1394 N$1393 "Straight Waveguide" sch_x=-59 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W698 N$1396 N$1395 "Straight Waveguide" sch_x=-59 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W699 N$1398 N$1397 "Straight Waveguide" sch_x=-57 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W700 N$1400 N$1399 "Straight Waveguide" sch_x=-57 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W701 N$1402 N$1401 "Straight Waveguide" sch_x=-57 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W702 N$1404 N$1403 "Straight Waveguide" sch_x=-57 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W703 N$1406 N$1405 "Straight Waveguide" sch_x=-57 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W704 N$1408 N$1407 "Straight Waveguide" sch_x=-57 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W705 N$1410 N$1409 "Straight Waveguide" sch_x=-57 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W706 N$1412 N$1411 "Straight Waveguide" sch_x=-57 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W707 N$1414 N$1413 "Straight Waveguide" sch_x=-57 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W708 N$1416 N$1415 "Straight Waveguide" sch_x=-57 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W709 N$1418 N$1417 "Straight Waveguide" sch_x=-57 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W710 N$1420 N$1419 "Straight Waveguide" sch_x=-57 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W711 N$1422 N$1421 "Straight Waveguide" sch_x=-57 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W712 N$1424 N$1423 "Straight Waveguide" sch_x=-57 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W713 N$1426 N$1425 "Straight Waveguide" sch_x=-57 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W714 N$1428 N$1427 "Straight Waveguide" sch_x=-57 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W715 N$1430 N$1429 "Straight Waveguide" sch_x=-57 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W716 N$1432 N$1431 "Straight Waveguide" sch_x=-57 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W717 N$1434 N$1433 "Straight Waveguide" sch_x=-57 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W718 N$1436 N$1435 "Straight Waveguide" sch_x=-57 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W719 N$1438 N$1437 "Straight Waveguide" sch_x=-57 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W720 N$1440 N$1439 "Straight Waveguide" sch_x=-57 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W721 N$1442 N$1441 "Straight Waveguide" sch_x=-57 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W722 N$1444 N$1443 "Straight Waveguide" sch_x=-57 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W723 N$1446 N$1445 "Straight Waveguide" sch_x=-57 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W724 N$1448 N$1447 "Straight Waveguide" sch_x=-57 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W725 N$1450 N$1449 "Straight Waveguide" sch_x=-55 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W726 N$1452 N$1451 "Straight Waveguide" sch_x=-55 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W727 N$1454 N$1453 "Straight Waveguide" sch_x=-55 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W728 N$1456 N$1455 "Straight Waveguide" sch_x=-55 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W729 N$1458 N$1457 "Straight Waveguide" sch_x=-55 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W730 N$1460 N$1459 "Straight Waveguide" sch_x=-55 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W731 N$1462 N$1461 "Straight Waveguide" sch_x=-55 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W732 N$1464 N$1463 "Straight Waveguide" sch_x=-55 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W733 N$1466 N$1465 "Straight Waveguide" sch_x=-55 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W734 N$1468 N$1467 "Straight Waveguide" sch_x=-55 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W735 N$1470 N$1469 "Straight Waveguide" sch_x=-55 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W736 N$1472 N$1471 "Straight Waveguide" sch_x=-55 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W737 N$1474 N$1473 "Straight Waveguide" sch_x=-55 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W738 N$1476 N$1475 "Straight Waveguide" sch_x=-55 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W739 N$1478 N$1477 "Straight Waveguide" sch_x=-55 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W740 N$1480 N$1479 "Straight Waveguide" sch_x=-55 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W741 N$1482 N$1481 "Straight Waveguide" sch_x=-55 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W742 N$1484 N$1483 "Straight Waveguide" sch_x=-55 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W743 N$1486 N$1485 "Straight Waveguide" sch_x=-55 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W744 N$1488 N$1487 "Straight Waveguide" sch_x=-55 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W745 N$1490 N$1489 "Straight Waveguide" sch_x=-55 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W746 N$1492 N$1491 "Straight Waveguide" sch_x=-55 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W747 N$1494 N$1493 "Straight Waveguide" sch_x=-55 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W748 N$1496 N$1495 "Straight Waveguide" sch_x=-55 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W749 N$1498 N$1497 "Straight Waveguide" sch_x=-53 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W750 N$1500 N$1499 "Straight Waveguide" sch_x=-53 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W751 N$1502 N$1501 "Straight Waveguide" sch_x=-53 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W752 N$1504 N$1503 "Straight Waveguide" sch_x=-53 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W753 N$1506 N$1505 "Straight Waveguide" sch_x=-53 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W754 N$1508 N$1507 "Straight Waveguide" sch_x=-53 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W755 N$1510 N$1509 "Straight Waveguide" sch_x=-53 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W756 N$1512 N$1511 "Straight Waveguide" sch_x=-53 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W757 N$1514 N$1513 "Straight Waveguide" sch_x=-53 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W758 N$1516 N$1515 "Straight Waveguide" sch_x=-53 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W759 N$1518 N$1517 "Straight Waveguide" sch_x=-53 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W760 N$1520 N$1519 "Straight Waveguide" sch_x=-53 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W761 N$1522 N$1521 "Straight Waveguide" sch_x=-53 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W762 N$1524 N$1523 "Straight Waveguide" sch_x=-53 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W763 N$1526 N$1525 "Straight Waveguide" sch_x=-53 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W764 N$1528 N$1527 "Straight Waveguide" sch_x=-53 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W765 N$1530 N$1529 "Straight Waveguide" sch_x=-53 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W766 N$1532 N$1531 "Straight Waveguide" sch_x=-53 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W767 N$1534 N$1533 "Straight Waveguide" sch_x=-53 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W768 N$1536 N$1535 "Straight Waveguide" sch_x=-53 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W769 N$1538 N$1537 "Straight Waveguide" sch_x=-53 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W770 N$1540 N$1539 "Straight Waveguide" sch_x=-53 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W771 N$1542 N$1541 "Straight Waveguide" sch_x=-51 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W772 N$1544 N$1543 "Straight Waveguide" sch_x=-51 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W773 N$1546 N$1545 "Straight Waveguide" sch_x=-51 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W774 N$1548 N$1547 "Straight Waveguide" sch_x=-51 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W775 N$1550 N$1549 "Straight Waveguide" sch_x=-51 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W776 N$1552 N$1551 "Straight Waveguide" sch_x=-51 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W777 N$1554 N$1553 "Straight Waveguide" sch_x=-51 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W778 N$1556 N$1555 "Straight Waveguide" sch_x=-51 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W779 N$1558 N$1557 "Straight Waveguide" sch_x=-51 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W780 N$1560 N$1559 "Straight Waveguide" sch_x=-51 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W781 N$1562 N$1561 "Straight Waveguide" sch_x=-51 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W782 N$1564 N$1563 "Straight Waveguide" sch_x=-51 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W783 N$1566 N$1565 "Straight Waveguide" sch_x=-51 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W784 N$1568 N$1567 "Straight Waveguide" sch_x=-51 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W785 N$1570 N$1569 "Straight Waveguide" sch_x=-51 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W786 N$1572 N$1571 "Straight Waveguide" sch_x=-51 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W787 N$1574 N$1573 "Straight Waveguide" sch_x=-51 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W788 N$1576 N$1575 "Straight Waveguide" sch_x=-51 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W789 N$1578 N$1577 "Straight Waveguide" sch_x=-51 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W790 N$1580 N$1579 "Straight Waveguide" sch_x=-51 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W791 N$1582 N$1581 "Straight Waveguide" sch_x=-49 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W792 N$1584 N$1583 "Straight Waveguide" sch_x=-49 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W793 N$1586 N$1585 "Straight Waveguide" sch_x=-49 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W794 N$1588 N$1587 "Straight Waveguide" sch_x=-49 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W795 N$1590 N$1589 "Straight Waveguide" sch_x=-49 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W796 N$1592 N$1591 "Straight Waveguide" sch_x=-49 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W797 N$1594 N$1593 "Straight Waveguide" sch_x=-49 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W798 N$1596 N$1595 "Straight Waveguide" sch_x=-49 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W799 N$1598 N$1597 "Straight Waveguide" sch_x=-49 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W800 N$1600 N$1599 "Straight Waveguide" sch_x=-49 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W801 N$1602 N$1601 "Straight Waveguide" sch_x=-49 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W802 N$1604 N$1603 "Straight Waveguide" sch_x=-49 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W803 N$1606 N$1605 "Straight Waveguide" sch_x=-49 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W804 N$1608 N$1607 "Straight Waveguide" sch_x=-49 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W805 N$1610 N$1609 "Straight Waveguide" sch_x=-49 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W806 N$1612 N$1611 "Straight Waveguide" sch_x=-49 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W807 N$1614 N$1613 "Straight Waveguide" sch_x=-49 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W808 N$1616 N$1615 "Straight Waveguide" sch_x=-49 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W809 N$1618 N$1617 "Straight Waveguide" sch_x=-47 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W810 N$1620 N$1619 "Straight Waveguide" sch_x=-47 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W811 N$1622 N$1621 "Straight Waveguide" sch_x=-47 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W812 N$1624 N$1623 "Straight Waveguide" sch_x=-47 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W813 N$1626 N$1625 "Straight Waveguide" sch_x=-47 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W814 N$1628 N$1627 "Straight Waveguide" sch_x=-47 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W815 N$1630 N$1629 "Straight Waveguide" sch_x=-47 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W816 N$1632 N$1631 "Straight Waveguide" sch_x=-47 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W817 N$1634 N$1633 "Straight Waveguide" sch_x=-47 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W818 N$1636 N$1635 "Straight Waveguide" sch_x=-47 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W819 N$1638 N$1637 "Straight Waveguide" sch_x=-47 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W820 N$1640 N$1639 "Straight Waveguide" sch_x=-47 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W821 N$1642 N$1641 "Straight Waveguide" sch_x=-47 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W822 N$1644 N$1643 "Straight Waveguide" sch_x=-47 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W823 N$1646 N$1645 "Straight Waveguide" sch_x=-47 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W824 N$1648 N$1647 "Straight Waveguide" sch_x=-47 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W825 N$1650 N$1649 "Straight Waveguide" sch_x=-45 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W826 N$1652 N$1651 "Straight Waveguide" sch_x=-45 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W827 N$1654 N$1653 "Straight Waveguide" sch_x=-45 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W828 N$1656 N$1655 "Straight Waveguide" sch_x=-45 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W829 N$1658 N$1657 "Straight Waveguide" sch_x=-45 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W830 N$1660 N$1659 "Straight Waveguide" sch_x=-45 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W831 N$1662 N$1661 "Straight Waveguide" sch_x=-45 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W832 N$1664 N$1663 "Straight Waveguide" sch_x=-45 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W833 N$1666 N$1665 "Straight Waveguide" sch_x=-45 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W834 N$1668 N$1667 "Straight Waveguide" sch_x=-45 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W835 N$1670 N$1669 "Straight Waveguide" sch_x=-45 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W836 N$1672 N$1671 "Straight Waveguide" sch_x=-45 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W837 N$1674 N$1673 "Straight Waveguide" sch_x=-45 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W838 N$1676 N$1675 "Straight Waveguide" sch_x=-45 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W839 N$1678 N$1677 "Straight Waveguide" sch_x=-43 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W840 N$1680 N$1679 "Straight Waveguide" sch_x=-43 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W841 N$1682 N$1681 "Straight Waveguide" sch_x=-43 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W842 N$1684 N$1683 "Straight Waveguide" sch_x=-43 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W843 N$1686 N$1685 "Straight Waveguide" sch_x=-43 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W844 N$1688 N$1687 "Straight Waveguide" sch_x=-43 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W845 N$1690 N$1689 "Straight Waveguide" sch_x=-43 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W846 N$1692 N$1691 "Straight Waveguide" sch_x=-43 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W847 N$1694 N$1693 "Straight Waveguide" sch_x=-43 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W848 N$1696 N$1695 "Straight Waveguide" sch_x=-43 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W849 N$1698 N$1697 "Straight Waveguide" sch_x=-43 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W850 N$1700 N$1699 "Straight Waveguide" sch_x=-43 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W851 N$1702 N$1701 "Straight Waveguide" sch_x=-41 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W852 N$1704 N$1703 "Straight Waveguide" sch_x=-41 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W853 N$1706 N$1705 "Straight Waveguide" sch_x=-41 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W854 N$1708 N$1707 "Straight Waveguide" sch_x=-41 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W855 N$1710 N$1709 "Straight Waveguide" sch_x=-41 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W856 N$1712 N$1711 "Straight Waveguide" sch_x=-41 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W857 N$1714 N$1713 "Straight Waveguide" sch_x=-41 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W858 N$1716 N$1715 "Straight Waveguide" sch_x=-41 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W859 N$1718 N$1717 "Straight Waveguide" sch_x=-41 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W860 N$1720 N$1719 "Straight Waveguide" sch_x=-41 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W861 N$1722 N$1721 "Straight Waveguide" sch_x=-39 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W862 N$1724 N$1723 "Straight Waveguide" sch_x=-39 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W863 N$1726 N$1725 "Straight Waveguide" sch_x=-39 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W864 N$1728 N$1727 "Straight Waveguide" sch_x=-39 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W865 N$1730 N$1729 "Straight Waveguide" sch_x=-39 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W866 N$1732 N$1731 "Straight Waveguide" sch_x=-39 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W867 N$1734 N$1733 "Straight Waveguide" sch_x=-39 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W868 N$1736 N$1735 "Straight Waveguide" sch_x=-39 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W869 N$1738 N$1737 "Straight Waveguide" sch_x=-37 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W870 N$1740 N$1739 "Straight Waveguide" sch_x=-37 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W871 N$1742 N$1741 "Straight Waveguide" sch_x=-37 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W872 N$1744 N$1743 "Straight Waveguide" sch_x=-37 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W873 N$1746 N$1745 "Straight Waveguide" sch_x=-37 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W874 N$1748 N$1747 "Straight Waveguide" sch_x=-37 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W875 N$1750 N$1749 "Straight Waveguide" sch_x=-35 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W876 N$1752 N$1751 "Straight Waveguide" sch_x=-35 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W877 N$1754 N$1753 "Straight Waveguide" sch_x=-35 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W878 N$1756 N$1755 "Straight Waveguide" sch_x=-35 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W879 N$1758 N$1757 "Straight Waveguide" sch_x=-33 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W880 N$1760 N$1759 "Straight Waveguide" sch_x=-33 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W881 N$1761 N$1762 "Straight Waveguide" sch_x=-45 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W882 N$1763 N$1764 "Straight Waveguide" sch_x=-44 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W883 N$1765 N$1766 "Straight Waveguide" sch_x=-43 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W884 N$1767 N$1768 "Straight Waveguide" sch_x=-42 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W885 N$1769 N$1770 "Straight Waveguide" sch_x=-41 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W886 N$1771 N$1772 "Straight Waveguide" sch_x=-40 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W887 N$1773 N$1774 "Straight Waveguide" sch_x=-39 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W888 N$1775 N$1776 "Straight Waveguide" sch_x=-38 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W889 N$1777 N$1778 "Straight Waveguide" sch_x=-37 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W890 N$1779 N$1780 "Straight Waveguide" sch_x=-36 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W891 N$1781 N$1782 "Straight Waveguide" sch_x=-35 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W892 N$1783 N$1784 "Straight Waveguide" sch_x=-34 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W893 N$1785 N$1786 "Straight Waveguide" sch_x=-33 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W894 N$1787 N$1788 "Straight Waveguide" sch_x=-32 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W895 N$1789 N$1790 "Straight Waveguide" sch_x=-31 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W896 N$1791 N$1792 "Straight Waveguide" sch_x=-31 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W897 N$1793 N$1794 "Straight Waveguide" sch_x=-32 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W898 N$1795 N$1796 "Straight Waveguide" sch_x=-33 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W899 N$1797 N$1798 "Straight Waveguide" sch_x=-34 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W900 N$1799 N$1800 "Straight Waveguide" sch_x=-35 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W901 N$1801 N$1802 "Straight Waveguide" sch_x=-36 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W902 N$1803 N$1804 "Straight Waveguide" sch_x=-37 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W903 N$1805 N$1806 "Straight Waveguide" sch_x=-38 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W904 N$1807 N$1808 "Straight Waveguide" sch_x=-39 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W905 N$1809 N$1810 "Straight Waveguide" sch_x=-40 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W906 N$1811 N$1812 "Straight Waveguide" sch_x=-41 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W907 N$1813 N$1814 "Straight Waveguide" sch_x=-42 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W908 N$1815 N$1816 "Straight Waveguide" sch_x=-43 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W909 N$1817 N$1818 "Straight Waveguide" sch_x=-44 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W910 N$1819 N$1820 "Straight Waveguide" sch_x=-45 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W911 N$1821 N$1822 "Straight Waveguide" sch_x=-46 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W912 N$1823 N$1824 "Straight Waveguide" sch_x=-46 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W913 N$1825 N$1826 "Straight Waveguide" sch_x=61 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W914 N$1827 N$1828 "Straight Waveguide" sch_x=61 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W915 N$1829 N$1830 "Straight Waveguide" sch_x=61 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W916 N$1831 N$1832 "Straight Waveguide" sch_x=61 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W917 N$1833 N$1834 "Straight Waveguide" sch_x=61 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W918 N$1835 N$1836 "Straight Waveguide" sch_x=61 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W919 N$1837 N$1838 "Straight Waveguide" sch_x=61 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W920 N$1839 N$1840 "Straight Waveguide" sch_x=61 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W921 N$1841 N$1842 "Straight Waveguide" sch_x=61 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W922 N$1843 N$1844 "Straight Waveguide" sch_x=61 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W923 N$1845 N$1846 "Straight Waveguide" sch_x=61 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W924 N$1847 N$1848 "Straight Waveguide" sch_x=61 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W925 N$1849 N$1850 "Straight Waveguide" sch_x=61 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W926 N$1851 N$1852 "Straight Waveguide" sch_x=61 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W927 N$1853 N$1854 "Straight Waveguide" sch_x=61 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W928 N$1855 N$1856 "Straight Waveguide" sch_x=61 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W929 N$1857 N$1858 "Straight Waveguide" sch_x=61 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W930 N$1859 N$1860 "Straight Waveguide" sch_x=61 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W931 N$1861 N$1862 "Straight Waveguide" sch_x=61 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W932 N$1863 N$1864 "Straight Waveguide" sch_x=61 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W933 N$1865 N$1866 "Straight Waveguide" sch_x=61 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W934 N$1867 N$1868 "Straight Waveguide" sch_x=61 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W935 N$1869 N$1870 "Straight Waveguide" sch_x=61 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W936 N$1871 N$1872 "Straight Waveguide" sch_x=61 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W937 N$1873 N$1874 "Straight Waveguide" sch_x=61 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W938 N$1875 N$1876 "Straight Waveguide" sch_x=61 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W939 N$1877 N$1878 "Straight Waveguide" sch_x=61 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W940 N$1879 N$1880 "Straight Waveguide" sch_x=61 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W941 N$1881 N$1882 "Straight Waveguide" sch_x=61 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W942 N$1883 N$1884 "Straight Waveguide" sch_x=61 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W943 N$1885 N$1886 "Straight Waveguide" sch_x=59 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W944 N$1887 N$1888 "Straight Waveguide" sch_x=59 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W945 N$1889 N$1890 "Straight Waveguide" sch_x=59 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W946 N$1891 N$1892 "Straight Waveguide" sch_x=59 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W947 N$1893 N$1894 "Straight Waveguide" sch_x=59 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W948 N$1895 N$1896 "Straight Waveguide" sch_x=59 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W949 N$1897 N$1898 "Straight Waveguide" sch_x=59 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W950 N$1899 N$1900 "Straight Waveguide" sch_x=59 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W951 N$1901 N$1902 "Straight Waveguide" sch_x=59 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W952 N$1903 N$1904 "Straight Waveguide" sch_x=59 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W953 N$1905 N$1906 "Straight Waveguide" sch_x=59 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W954 N$1907 N$1908 "Straight Waveguide" sch_x=59 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W955 N$1909 N$1910 "Straight Waveguide" sch_x=59 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W956 N$1911 N$1912 "Straight Waveguide" sch_x=59 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W957 N$1913 N$1914 "Straight Waveguide" sch_x=59 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W958 N$1915 N$1916 "Straight Waveguide" sch_x=59 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W959 N$1917 N$1918 "Straight Waveguide" sch_x=59 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W960 N$1919 N$1920 "Straight Waveguide" sch_x=59 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W961 N$1921 N$1922 "Straight Waveguide" sch_x=59 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W962 N$1923 N$1924 "Straight Waveguide" sch_x=59 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W963 N$1925 N$1926 "Straight Waveguide" sch_x=59 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W964 N$1927 N$1928 "Straight Waveguide" sch_x=59 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W965 N$1929 N$1930 "Straight Waveguide" sch_x=59 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W966 N$1931 N$1932 "Straight Waveguide" sch_x=59 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W967 N$1933 N$1934 "Straight Waveguide" sch_x=59 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W968 N$1935 N$1936 "Straight Waveguide" sch_x=59 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W969 N$1937 N$1938 "Straight Waveguide" sch_x=59 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W970 N$1939 N$1940 "Straight Waveguide" sch_x=59 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W971 N$1941 N$1942 "Straight Waveguide" sch_x=57 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W972 N$1943 N$1944 "Straight Waveguide" sch_x=57 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W973 N$1945 N$1946 "Straight Waveguide" sch_x=57 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W974 N$1947 N$1948 "Straight Waveguide" sch_x=57 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W975 N$1949 N$1950 "Straight Waveguide" sch_x=57 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W976 N$1951 N$1952 "Straight Waveguide" sch_x=57 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W977 N$1953 N$1954 "Straight Waveguide" sch_x=57 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W978 N$1955 N$1956 "Straight Waveguide" sch_x=57 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W979 N$1957 N$1958 "Straight Waveguide" sch_x=57 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W980 N$1959 N$1960 "Straight Waveguide" sch_x=57 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W981 N$1961 N$1962 "Straight Waveguide" sch_x=57 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W982 N$1963 N$1964 "Straight Waveguide" sch_x=57 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W983 N$1965 N$1966 "Straight Waveguide" sch_x=57 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W984 N$1967 N$1968 "Straight Waveguide" sch_x=57 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W985 N$1969 N$1970 "Straight Waveguide" sch_x=57 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W986 N$1971 N$1972 "Straight Waveguide" sch_x=57 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W987 N$1973 N$1974 "Straight Waveguide" sch_x=57 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W988 N$1975 N$1976 "Straight Waveguide" sch_x=57 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W989 N$1977 N$1978 "Straight Waveguide" sch_x=57 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W990 N$1979 N$1980 "Straight Waveguide" sch_x=57 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W991 N$1981 N$1982 "Straight Waveguide" sch_x=57 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W992 N$1983 N$1984 "Straight Waveguide" sch_x=57 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W993 N$1985 N$1986 "Straight Waveguide" sch_x=57 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W994 N$1987 N$1988 "Straight Waveguide" sch_x=57 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W995 N$1989 N$1990 "Straight Waveguide" sch_x=57 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W996 N$1991 N$1992 "Straight Waveguide" sch_x=57 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W997 N$1993 N$1994 "Straight Waveguide" sch_x=55 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W998 N$1995 N$1996 "Straight Waveguide" sch_x=55 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W999 N$1997 N$1998 "Straight Waveguide" sch_x=55 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1000 N$1999 N$2000 "Straight Waveguide" sch_x=55 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1001 N$2001 N$2002 "Straight Waveguide" sch_x=55 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1002 N$2003 N$2004 "Straight Waveguide" sch_x=55 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1003 N$2005 N$2006 "Straight Waveguide" sch_x=55 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1004 N$2007 N$2008 "Straight Waveguide" sch_x=55 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1005 N$2009 N$2010 "Straight Waveguide" sch_x=55 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1006 N$2011 N$2012 "Straight Waveguide" sch_x=55 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1007 N$2013 N$2014 "Straight Waveguide" sch_x=55 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1008 N$2015 N$2016 "Straight Waveguide" sch_x=55 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1009 N$2017 N$2018 "Straight Waveguide" sch_x=55 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1010 N$2019 N$2020 "Straight Waveguide" sch_x=55 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1011 N$2021 N$2022 "Straight Waveguide" sch_x=55 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1012 N$2023 N$2024 "Straight Waveguide" sch_x=55 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1013 N$2025 N$2026 "Straight Waveguide" sch_x=55 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1014 N$2027 N$2028 "Straight Waveguide" sch_x=55 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1015 N$2029 N$2030 "Straight Waveguide" sch_x=55 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1016 N$2031 N$2032 "Straight Waveguide" sch_x=55 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1017 N$2033 N$2034 "Straight Waveguide" sch_x=55 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1018 N$2035 N$2036 "Straight Waveguide" sch_x=55 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1019 N$2037 N$2038 "Straight Waveguide" sch_x=55 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1020 N$2039 N$2040 "Straight Waveguide" sch_x=55 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1021 N$2041 N$2042 "Straight Waveguide" sch_x=53 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1022 N$2043 N$2044 "Straight Waveguide" sch_x=53 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1023 N$2045 N$2046 "Straight Waveguide" sch_x=53 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1024 N$2047 N$2048 "Straight Waveguide" sch_x=53 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1025 N$2049 N$2050 "Straight Waveguide" sch_x=53 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1026 N$2051 N$2052 "Straight Waveguide" sch_x=53 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1027 N$2053 N$2054 "Straight Waveguide" sch_x=53 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1028 N$2055 N$2056 "Straight Waveguide" sch_x=53 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1029 N$2057 N$2058 "Straight Waveguide" sch_x=53 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1030 N$2059 N$2060 "Straight Waveguide" sch_x=53 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1031 N$2061 N$2062 "Straight Waveguide" sch_x=53 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1032 N$2063 N$2064 "Straight Waveguide" sch_x=53 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1033 N$2065 N$2066 "Straight Waveguide" sch_x=53 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1034 N$2067 N$2068 "Straight Waveguide" sch_x=53 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1035 N$2069 N$2070 "Straight Waveguide" sch_x=53 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1036 N$2071 N$2072 "Straight Waveguide" sch_x=53 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1037 N$2073 N$2074 "Straight Waveguide" sch_x=53 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1038 N$2075 N$2076 "Straight Waveguide" sch_x=53 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1039 N$2077 N$2078 "Straight Waveguide" sch_x=53 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1040 N$2079 N$2080 "Straight Waveguide" sch_x=53 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1041 N$2081 N$2082 "Straight Waveguide" sch_x=53 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1042 N$2083 N$2084 "Straight Waveguide" sch_x=53 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1043 N$2085 N$2086 "Straight Waveguide" sch_x=51 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1044 N$2087 N$2088 "Straight Waveguide" sch_x=51 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1045 N$2089 N$2090 "Straight Waveguide" sch_x=51 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1046 N$2091 N$2092 "Straight Waveguide" sch_x=51 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1047 N$2093 N$2094 "Straight Waveguide" sch_x=51 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1048 N$2095 N$2096 "Straight Waveguide" sch_x=51 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1049 N$2097 N$2098 "Straight Waveguide" sch_x=51 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1050 N$2099 N$2100 "Straight Waveguide" sch_x=51 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1051 N$2101 N$2102 "Straight Waveguide" sch_x=51 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1052 N$2103 N$2104 "Straight Waveguide" sch_x=51 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1053 N$2105 N$2106 "Straight Waveguide" sch_x=51 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1054 N$2107 N$2108 "Straight Waveguide" sch_x=51 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1055 N$2109 N$2110 "Straight Waveguide" sch_x=51 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1056 N$2111 N$2112 "Straight Waveguide" sch_x=51 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1057 N$2113 N$2114 "Straight Waveguide" sch_x=51 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1058 N$2115 N$2116 "Straight Waveguide" sch_x=51 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1059 N$2117 N$2118 "Straight Waveguide" sch_x=51 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1060 N$2119 N$2120 "Straight Waveguide" sch_x=51 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1061 N$2121 N$2122 "Straight Waveguide" sch_x=51 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1062 N$2123 N$2124 "Straight Waveguide" sch_x=51 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1063 N$2125 N$2126 "Straight Waveguide" sch_x=49 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1064 N$2127 N$2128 "Straight Waveguide" sch_x=49 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1065 N$2129 N$2130 "Straight Waveguide" sch_x=49 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1066 N$2131 N$2132 "Straight Waveguide" sch_x=49 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1067 N$2133 N$2134 "Straight Waveguide" sch_x=49 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1068 N$2135 N$2136 "Straight Waveguide" sch_x=49 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1069 N$2137 N$2138 "Straight Waveguide" sch_x=49 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1070 N$2139 N$2140 "Straight Waveguide" sch_x=49 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1071 N$2141 N$2142 "Straight Waveguide" sch_x=49 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1072 N$2143 N$2144 "Straight Waveguide" sch_x=49 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1073 N$2145 N$2146 "Straight Waveguide" sch_x=49 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1074 N$2147 N$2148 "Straight Waveguide" sch_x=49 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1075 N$2149 N$2150 "Straight Waveguide" sch_x=49 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1076 N$2151 N$2152 "Straight Waveguide" sch_x=49 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1077 N$2153 N$2154 "Straight Waveguide" sch_x=49 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1078 N$2155 N$2156 "Straight Waveguide" sch_x=49 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1079 N$2157 N$2158 "Straight Waveguide" sch_x=49 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1080 N$2159 N$2160 "Straight Waveguide" sch_x=49 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1081 N$2161 N$2162 "Straight Waveguide" sch_x=47 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1082 N$2163 N$2164 "Straight Waveguide" sch_x=47 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1083 N$2165 N$2166 "Straight Waveguide" sch_x=47 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1084 N$2167 N$2168 "Straight Waveguide" sch_x=47 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1085 N$2169 N$2170 "Straight Waveguide" sch_x=47 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1086 N$2171 N$2172 "Straight Waveguide" sch_x=47 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1087 N$2173 N$2174 "Straight Waveguide" sch_x=47 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1088 N$2175 N$2176 "Straight Waveguide" sch_x=47 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1089 N$2177 N$2178 "Straight Waveguide" sch_x=47 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1090 N$2179 N$2180 "Straight Waveguide" sch_x=47 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1091 N$2181 N$2182 "Straight Waveguide" sch_x=47 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1092 N$2183 N$2184 "Straight Waveguide" sch_x=47 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1093 N$2185 N$2186 "Straight Waveguide" sch_x=47 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1094 N$2187 N$2188 "Straight Waveguide" sch_x=47 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1095 N$2189 N$2190 "Straight Waveguide" sch_x=47 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1096 N$2191 N$2192 "Straight Waveguide" sch_x=47 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1097 N$2193 N$2194 "Straight Waveguide" sch_x=45 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1098 N$2195 N$2196 "Straight Waveguide" sch_x=45 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1099 N$2197 N$2198 "Straight Waveguide" sch_x=45 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1100 N$2199 N$2200 "Straight Waveguide" sch_x=45 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1101 N$2201 N$2202 "Straight Waveguide" sch_x=45 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1102 N$2203 N$2204 "Straight Waveguide" sch_x=45 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1103 N$2205 N$2206 "Straight Waveguide" sch_x=45 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1104 N$2207 N$2208 "Straight Waveguide" sch_x=45 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1105 N$2209 N$2210 "Straight Waveguide" sch_x=45 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1106 N$2211 N$2212 "Straight Waveguide" sch_x=45 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1107 N$2213 N$2214 "Straight Waveguide" sch_x=45 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1108 N$2215 N$2216 "Straight Waveguide" sch_x=45 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1109 N$2217 N$2218 "Straight Waveguide" sch_x=45 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1110 N$2219 N$2220 "Straight Waveguide" sch_x=45 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1111 N$2221 N$2222 "Straight Waveguide" sch_x=43 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1112 N$2223 N$2224 "Straight Waveguide" sch_x=43 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1113 N$2225 N$2226 "Straight Waveguide" sch_x=43 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1114 N$2227 N$2228 "Straight Waveguide" sch_x=43 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1115 N$2229 N$2230 "Straight Waveguide" sch_x=43 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1116 N$2231 N$2232 "Straight Waveguide" sch_x=43 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1117 N$2233 N$2234 "Straight Waveguide" sch_x=43 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1118 N$2235 N$2236 "Straight Waveguide" sch_x=43 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1119 N$2237 N$2238 "Straight Waveguide" sch_x=43 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1120 N$2239 N$2240 "Straight Waveguide" sch_x=43 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1121 N$2241 N$2242 "Straight Waveguide" sch_x=43 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1122 N$2243 N$2244 "Straight Waveguide" sch_x=43 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1123 N$2245 N$2246 "Straight Waveguide" sch_x=41 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1124 N$2247 N$2248 "Straight Waveguide" sch_x=41 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1125 N$2249 N$2250 "Straight Waveguide" sch_x=41 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1126 N$2251 N$2252 "Straight Waveguide" sch_x=41 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1127 N$2253 N$2254 "Straight Waveguide" sch_x=41 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1128 N$2255 N$2256 "Straight Waveguide" sch_x=41 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1129 N$2257 N$2258 "Straight Waveguide" sch_x=41 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1130 N$2259 N$2260 "Straight Waveguide" sch_x=41 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1131 N$2261 N$2262 "Straight Waveguide" sch_x=41 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1132 N$2263 N$2264 "Straight Waveguide" sch_x=41 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1133 N$2265 N$2266 "Straight Waveguide" sch_x=39 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1134 N$2267 N$2268 "Straight Waveguide" sch_x=39 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1135 N$2269 N$2270 "Straight Waveguide" sch_x=39 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1136 N$2271 N$2272 "Straight Waveguide" sch_x=39 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1137 N$2273 N$2274 "Straight Waveguide" sch_x=39 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1138 N$2275 N$2276 "Straight Waveguide" sch_x=39 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1139 N$2277 N$2278 "Straight Waveguide" sch_x=39 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1140 N$2279 N$2280 "Straight Waveguide" sch_x=39 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1141 N$2281 N$2282 "Straight Waveguide" sch_x=37 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1142 N$2283 N$2284 "Straight Waveguide" sch_x=37 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1143 N$2285 N$2286 "Straight Waveguide" sch_x=37 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1144 N$2287 N$2288 "Straight Waveguide" sch_x=37 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1145 N$2289 N$2290 "Straight Waveguide" sch_x=37 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1146 N$2291 N$2292 "Straight Waveguide" sch_x=37 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1147 N$2293 N$2294 "Straight Waveguide" sch_x=35 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1148 N$2295 N$2296 "Straight Waveguide" sch_x=35 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1149 N$2297 N$2298 "Straight Waveguide" sch_x=35 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1150 N$2299 N$2300 "Straight Waveguide" sch_x=35 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1151 N$2301 N$2302 "Straight Waveguide" sch_x=33 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1152 N$2303 N$2304 "Straight Waveguide" sch_x=33 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1153 N$2306 N$2305 "Straight Waveguide" sch_x=45 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1154 N$2308 N$2307 "Straight Waveguide" sch_x=44 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1155 N$2310 N$2309 "Straight Waveguide" sch_x=43 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1156 N$2312 N$2311 "Straight Waveguide" sch_x=42 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1157 N$2314 N$2313 "Straight Waveguide" sch_x=41 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1158 N$2316 N$2315 "Straight Waveguide" sch_x=40 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1159 N$2318 N$2317 "Straight Waveguide" sch_x=39 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1160 N$2320 N$2319 "Straight Waveguide" sch_x=38 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1161 N$2322 N$2321 "Straight Waveguide" sch_x=37 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1162 N$2324 N$2323 "Straight Waveguide" sch_x=36 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1163 N$2326 N$2325 "Straight Waveguide" sch_x=35 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1164 N$2328 N$2327 "Straight Waveguide" sch_x=34 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1165 N$2330 N$2329 "Straight Waveguide" sch_x=33 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1166 N$2332 N$2331 "Straight Waveguide" sch_x=32 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1167 N$2334 N$2333 "Straight Waveguide" sch_x=31 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1168 N$2336 N$2335 "Straight Waveguide" sch_x=31 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1169 N$2338 N$2337 "Straight Waveguide" sch_x=32 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1170 N$2340 N$2339 "Straight Waveguide" sch_x=33 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1171 N$2342 N$2341 "Straight Waveguide" sch_x=34 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1172 N$2344 N$2343 "Straight Waveguide" sch_x=35 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1173 N$2346 N$2345 "Straight Waveguide" sch_x=36 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1174 N$2348 N$2347 "Straight Waveguide" sch_x=37 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1175 N$2350 N$2349 "Straight Waveguide" sch_x=38 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1176 N$2352 N$2351 "Straight Waveguide" sch_x=39 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1177 N$2354 N$2353 "Straight Waveguide" sch_x=40 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1178 N$2356 N$2355 "Straight Waveguide" sch_x=41 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1179 N$2358 N$2357 "Straight Waveguide" sch_x=42 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1180 N$2360 N$2359 "Straight Waveguide" sch_x=43 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1181 N$2362 N$2361 "Straight Waveguide" sch_x=44 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1182 N$2364 N$2363 "Straight Waveguide" sch_x=45 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1183 N$2366 N$2365 "Straight Waveguide" sch_x=46 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1184 N$2368 N$2367 "Straight Waveguide" sch_x=46 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1185 N$2369 N$2370 "Straight Waveguide" sch_x=-4 sch_y=31.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1186 N$2371 N$2372 "Straight Waveguide" sch_x=-5 sch_y=30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1187 N$2373 N$2374 "Straight Waveguide" sch_x=-5 sch_y=29.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1188 N$2375 N$2376 "Straight Waveguide" sch_x=-3 sch_y=30.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1189 N$2377 N$2378 "Straight Waveguide" sch_x=-3 sch_y=29.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1190 N$2379 N$2380 "Straight Waveguide" sch_x=-4 sch_y=28.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1191 N$2381 N$2382 "Straight Waveguide" sch_x=0 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1192 N$2383 N$2384 "Straight Waveguide" sch_x=-1 sch_y=31.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1193 N$2385 N$2386 "Straight Waveguide" sch_x=-1 sch_y=30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1194 N$2387 N$2388 "Straight Waveguide" sch_x=1 sch_y=30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1195 N$2389 N$2390 "Straight Waveguide" sch_x=1 sch_y=31.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1196 N$2391 N$2392 "Straight Waveguide" sch_x=0 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1197 N$2393 N$2394 "Straight Waveguide" sch_x=0 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1198 N$2395 N$2396 "Straight Waveguide" sch_x=-1 sch_y=29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1199 N$2397 N$2398 "Straight Waveguide" sch_x=-1 sch_y=28.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1200 N$2399 N$2400 "Straight Waveguide" sch_x=1 sch_y=28.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1201 N$2401 N$2402 "Straight Waveguide" sch_x=1 sch_y=29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1202 N$2403 N$2404 "Straight Waveguide" sch_x=0 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1203 N$2405 N$2406 "Straight Waveguide" sch_x=4 sch_y=31.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1204 N$2407 N$2408 "Straight Waveguide" sch_x=3 sch_y=30.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1205 N$2409 N$2410 "Straight Waveguide" sch_x=3 sch_y=29.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1206 N$2411 N$2412 "Straight Waveguide" sch_x=5 sch_y=29.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1207 N$2413 N$2414 "Straight Waveguide" sch_x=5 sch_y=30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1208 N$2415 N$2416 "Straight Waveguide" sch_x=4 sch_y=28.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1209 N$2417 N$2418 "Straight Waveguide" sch_x=-4 sch_y=27.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1210 N$2419 N$2420 "Straight Waveguide" sch_x=-5 sch_y=26.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1211 N$2421 N$2422 "Straight Waveguide" sch_x=-5 sch_y=25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1212 N$2423 N$2424 "Straight Waveguide" sch_x=-3 sch_y=26.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1213 N$2425 N$2426 "Straight Waveguide" sch_x=-3 sch_y=25.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1214 N$2427 N$2428 "Straight Waveguide" sch_x=-4 sch_y=24.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1215 N$2429 N$2430 "Straight Waveguide" sch_x=0 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1216 N$2431 N$2432 "Straight Waveguide" sch_x=-1 sch_y=27.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1217 N$2433 N$2434 "Straight Waveguide" sch_x=-1 sch_y=26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1218 N$2435 N$2436 "Straight Waveguide" sch_x=1 sch_y=26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1219 N$2437 N$2438 "Straight Waveguide" sch_x=1 sch_y=27.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1220 N$2439 N$2440 "Straight Waveguide" sch_x=0 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1221 N$2441 N$2442 "Straight Waveguide" sch_x=0 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1222 N$2443 N$2444 "Straight Waveguide" sch_x=-1 sch_y=25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1223 N$2445 N$2446 "Straight Waveguide" sch_x=-1 sch_y=24.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1224 N$2447 N$2448 "Straight Waveguide" sch_x=1 sch_y=24.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1225 N$2449 N$2450 "Straight Waveguide" sch_x=1 sch_y=25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1226 N$2451 N$2452 "Straight Waveguide" sch_x=0 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1227 N$2453 N$2454 "Straight Waveguide" sch_x=4 sch_y=27.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1228 N$2455 N$2456 "Straight Waveguide" sch_x=3 sch_y=26.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1229 N$2457 N$2458 "Straight Waveguide" sch_x=3 sch_y=25.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1230 N$2459 N$2460 "Straight Waveguide" sch_x=5 sch_y=25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1231 N$2461 N$2462 "Straight Waveguide" sch_x=5 sch_y=26.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1232 N$2463 N$2464 "Straight Waveguide" sch_x=4 sch_y=24.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1233 N$2466 N$2465 "Straight Waveguide" sch_x=-13 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1234 N$2468 N$2467 "Straight Waveguide" sch_x=-13 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1235 N$2470 N$2469 "Straight Waveguide" sch_x=-13 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1236 N$2472 N$2471 "Straight Waveguide" sch_x=-13 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1237 N$2474 N$2473 "Straight Waveguide" sch_x=-13 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1238 N$2476 N$2475 "Straight Waveguide" sch_x=-13 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1239 N$2478 N$2477 "Straight Waveguide" sch_x=-11 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1240 N$2480 N$2479 "Straight Waveguide" sch_x=-11 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1241 N$2482 N$2481 "Straight Waveguide" sch_x=-11 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1242 N$2484 N$2483 "Straight Waveguide" sch_x=-11 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1243 N$2486 N$2485 "Straight Waveguide" sch_x=-9 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1244 N$2488 N$2487 "Straight Waveguide" sch_x=-9 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1245 N$2489 N$2490 "Straight Waveguide" sch_x=-9 sch_y=30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1246 N$2491 N$2492 "Straight Waveguide" sch_x=-8 sch_y=29.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1247 N$2493 N$2494 "Straight Waveguide" sch_x=-7 sch_y=28.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1248 N$2495 N$2496 "Straight Waveguide" sch_x=-7 sch_y=27.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1249 N$2497 N$2498 "Straight Waveguide" sch_x=-8 sch_y=26.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1250 N$2499 N$2500 "Straight Waveguide" sch_x=-9 sch_y=25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1251 N$2501 N$2502 "Straight Waveguide" sch_x=-10 sch_y=30.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1252 N$2503 N$2504 "Straight Waveguide" sch_x=-10 sch_y=25.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1253 N$2505 N$2506 "Straight Waveguide" sch_x=13 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1254 N$2507 N$2508 "Straight Waveguide" sch_x=13 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1255 N$2509 N$2510 "Straight Waveguide" sch_x=13 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1256 N$2511 N$2512 "Straight Waveguide" sch_x=13 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1257 N$2513 N$2514 "Straight Waveguide" sch_x=13 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1258 N$2515 N$2516 "Straight Waveguide" sch_x=13 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1259 N$2517 N$2518 "Straight Waveguide" sch_x=11 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1260 N$2519 N$2520 "Straight Waveguide" sch_x=11 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1261 N$2521 N$2522 "Straight Waveguide" sch_x=11 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1262 N$2523 N$2524 "Straight Waveguide" sch_x=11 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1263 N$2525 N$2526 "Straight Waveguide" sch_x=9 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1264 N$2527 N$2528 "Straight Waveguide" sch_x=9 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1265 N$2530 N$2529 "Straight Waveguide" sch_x=9 sch_y=30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1266 N$2532 N$2531 "Straight Waveguide" sch_x=8 sch_y=29.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1267 N$2534 N$2533 "Straight Waveguide" sch_x=7 sch_y=28.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1268 N$2536 N$2535 "Straight Waveguide" sch_x=7 sch_y=27.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1269 N$2538 N$2537 "Straight Waveguide" sch_x=8 sch_y=26.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1270 N$2540 N$2539 "Straight Waveguide" sch_x=9 sch_y=25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1271 N$2542 N$2541 "Straight Waveguide" sch_x=10 sch_y=30.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1272 N$2544 N$2543 "Straight Waveguide" sch_x=10 sch_y=25.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1273 N$2545 N$2546 "Straight Waveguide" sch_x=-4 sch_y=23.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1274 N$2547 N$2548 "Straight Waveguide" sch_x=-5 sch_y=22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1275 N$2549 N$2550 "Straight Waveguide" sch_x=-5 sch_y=21.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1276 N$2551 N$2552 "Straight Waveguide" sch_x=-3 sch_y=22.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1277 N$2553 N$2554 "Straight Waveguide" sch_x=-3 sch_y=21.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1278 N$2555 N$2556 "Straight Waveguide" sch_x=-4 sch_y=20.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1279 N$2557 N$2558 "Straight Waveguide" sch_x=0 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1280 N$2559 N$2560 "Straight Waveguide" sch_x=-1 sch_y=23.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1281 N$2561 N$2562 "Straight Waveguide" sch_x=-1 sch_y=22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1282 N$2563 N$2564 "Straight Waveguide" sch_x=1 sch_y=22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1283 N$2565 N$2566 "Straight Waveguide" sch_x=1 sch_y=23.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1284 N$2567 N$2568 "Straight Waveguide" sch_x=0 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1285 N$2569 N$2570 "Straight Waveguide" sch_x=0 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1286 N$2571 N$2572 "Straight Waveguide" sch_x=-1 sch_y=21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1287 N$2573 N$2574 "Straight Waveguide" sch_x=-1 sch_y=20.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1288 N$2575 N$2576 "Straight Waveguide" sch_x=1 sch_y=20.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1289 N$2577 N$2578 "Straight Waveguide" sch_x=1 sch_y=21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1290 N$2579 N$2580 "Straight Waveguide" sch_x=0 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1291 N$2581 N$2582 "Straight Waveguide" sch_x=4 sch_y=23.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1292 N$2583 N$2584 "Straight Waveguide" sch_x=3 sch_y=22.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1293 N$2585 N$2586 "Straight Waveguide" sch_x=3 sch_y=21.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1294 N$2587 N$2588 "Straight Waveguide" sch_x=5 sch_y=21.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1295 N$2589 N$2590 "Straight Waveguide" sch_x=5 sch_y=22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1296 N$2591 N$2592 "Straight Waveguide" sch_x=4 sch_y=20.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1297 N$2593 N$2594 "Straight Waveguide" sch_x=-4 sch_y=19.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1298 N$2595 N$2596 "Straight Waveguide" sch_x=-5 sch_y=18.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1299 N$2597 N$2598 "Straight Waveguide" sch_x=-5 sch_y=17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1300 N$2599 N$2600 "Straight Waveguide" sch_x=-3 sch_y=18.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1301 N$2601 N$2602 "Straight Waveguide" sch_x=-3 sch_y=17.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1302 N$2603 N$2604 "Straight Waveguide" sch_x=-4 sch_y=16.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1303 N$2605 N$2606 "Straight Waveguide" sch_x=0 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1304 N$2607 N$2608 "Straight Waveguide" sch_x=-1 sch_y=19.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1305 N$2609 N$2610 "Straight Waveguide" sch_x=-1 sch_y=18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1306 N$2611 N$2612 "Straight Waveguide" sch_x=1 sch_y=18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1307 N$2613 N$2614 "Straight Waveguide" sch_x=1 sch_y=19.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1308 N$2615 N$2616 "Straight Waveguide" sch_x=0 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1309 N$2617 N$2618 "Straight Waveguide" sch_x=0 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1310 N$2619 N$2620 "Straight Waveguide" sch_x=-1 sch_y=17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1311 N$2621 N$2622 "Straight Waveguide" sch_x=-1 sch_y=16.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1312 N$2623 N$2624 "Straight Waveguide" sch_x=1 sch_y=16.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1313 N$2625 N$2626 "Straight Waveguide" sch_x=1 sch_y=17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1314 N$2627 N$2628 "Straight Waveguide" sch_x=0 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1315 N$2629 N$2630 "Straight Waveguide" sch_x=4 sch_y=19.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1316 N$2631 N$2632 "Straight Waveguide" sch_x=3 sch_y=18.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1317 N$2633 N$2634 "Straight Waveguide" sch_x=3 sch_y=17.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1318 N$2635 N$2636 "Straight Waveguide" sch_x=5 sch_y=17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1319 N$2637 N$2638 "Straight Waveguide" sch_x=5 sch_y=18.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1320 N$2639 N$2640 "Straight Waveguide" sch_x=4 sch_y=16.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1321 N$2642 N$2641 "Straight Waveguide" sch_x=-13 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1322 N$2644 N$2643 "Straight Waveguide" sch_x=-13 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1323 N$2646 N$2645 "Straight Waveguide" sch_x=-13 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1324 N$2648 N$2647 "Straight Waveguide" sch_x=-13 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1325 N$2650 N$2649 "Straight Waveguide" sch_x=-13 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1326 N$2652 N$2651 "Straight Waveguide" sch_x=-13 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1327 N$2654 N$2653 "Straight Waveguide" sch_x=-11 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1328 N$2656 N$2655 "Straight Waveguide" sch_x=-11 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1329 N$2658 N$2657 "Straight Waveguide" sch_x=-11 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1330 N$2660 N$2659 "Straight Waveguide" sch_x=-11 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1331 N$2662 N$2661 "Straight Waveguide" sch_x=-9 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1332 N$2664 N$2663 "Straight Waveguide" sch_x=-9 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1333 N$2665 N$2666 "Straight Waveguide" sch_x=-9 sch_y=22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1334 N$2667 N$2668 "Straight Waveguide" sch_x=-8 sch_y=21.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1335 N$2669 N$2670 "Straight Waveguide" sch_x=-7 sch_y=20.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1336 N$2671 N$2672 "Straight Waveguide" sch_x=-7 sch_y=19.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1337 N$2673 N$2674 "Straight Waveguide" sch_x=-8 sch_y=18.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1338 N$2675 N$2676 "Straight Waveguide" sch_x=-9 sch_y=17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1339 N$2677 N$2678 "Straight Waveguide" sch_x=-10 sch_y=22.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1340 N$2679 N$2680 "Straight Waveguide" sch_x=-10 sch_y=17.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1341 N$2681 N$2682 "Straight Waveguide" sch_x=13 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1342 N$2683 N$2684 "Straight Waveguide" sch_x=13 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1343 N$2685 N$2686 "Straight Waveguide" sch_x=13 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1344 N$2687 N$2688 "Straight Waveguide" sch_x=13 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1345 N$2689 N$2690 "Straight Waveguide" sch_x=13 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1346 N$2691 N$2692 "Straight Waveguide" sch_x=13 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1347 N$2693 N$2694 "Straight Waveguide" sch_x=11 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1348 N$2695 N$2696 "Straight Waveguide" sch_x=11 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1349 N$2697 N$2698 "Straight Waveguide" sch_x=11 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1350 N$2699 N$2700 "Straight Waveguide" sch_x=11 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1351 N$2701 N$2702 "Straight Waveguide" sch_x=9 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1352 N$2703 N$2704 "Straight Waveguide" sch_x=9 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1353 N$2706 N$2705 "Straight Waveguide" sch_x=9 sch_y=22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1354 N$2708 N$2707 "Straight Waveguide" sch_x=8 sch_y=21.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1355 N$2710 N$2709 "Straight Waveguide" sch_x=7 sch_y=20.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1356 N$2712 N$2711 "Straight Waveguide" sch_x=7 sch_y=19.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1357 N$2714 N$2713 "Straight Waveguide" sch_x=8 sch_y=18.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1358 N$2716 N$2715 "Straight Waveguide" sch_x=9 sch_y=17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1359 N$2718 N$2717 "Straight Waveguide" sch_x=10 sch_y=22.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1360 N$2720 N$2719 "Straight Waveguide" sch_x=10 sch_y=17.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1361 N$2722 N$2721 "Straight Waveguide" sch_x=-29 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1362 N$2724 N$2723 "Straight Waveguide" sch_x=-29 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1363 N$2726 N$2725 "Straight Waveguide" sch_x=-29 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1364 N$2728 N$2727 "Straight Waveguide" sch_x=-29 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1365 N$2730 N$2729 "Straight Waveguide" sch_x=-29 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1366 N$2732 N$2731 "Straight Waveguide" sch_x=-29 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1367 N$2734 N$2733 "Straight Waveguide" sch_x=-29 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1368 N$2736 N$2735 "Straight Waveguide" sch_x=-29 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1369 N$2738 N$2737 "Straight Waveguide" sch_x=-29 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1370 N$2740 N$2739 "Straight Waveguide" sch_x=-29 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1371 N$2742 N$2741 "Straight Waveguide" sch_x=-29 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1372 N$2744 N$2743 "Straight Waveguide" sch_x=-29 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1373 N$2746 N$2745 "Straight Waveguide" sch_x=-29 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1374 N$2748 N$2747 "Straight Waveguide" sch_x=-29 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1375 N$2750 N$2749 "Straight Waveguide" sch_x=-27 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1376 N$2752 N$2751 "Straight Waveguide" sch_x=-27 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1377 N$2754 N$2753 "Straight Waveguide" sch_x=-27 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1378 N$2756 N$2755 "Straight Waveguide" sch_x=-27 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1379 N$2758 N$2757 "Straight Waveguide" sch_x=-27 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1380 N$2760 N$2759 "Straight Waveguide" sch_x=-27 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1381 N$2762 N$2761 "Straight Waveguide" sch_x=-27 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1382 N$2764 N$2763 "Straight Waveguide" sch_x=-27 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1383 N$2766 N$2765 "Straight Waveguide" sch_x=-27 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1384 N$2768 N$2767 "Straight Waveguide" sch_x=-27 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1385 N$2770 N$2769 "Straight Waveguide" sch_x=-27 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1386 N$2772 N$2771 "Straight Waveguide" sch_x=-27 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1387 N$2774 N$2773 "Straight Waveguide" sch_x=-25 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1388 N$2776 N$2775 "Straight Waveguide" sch_x=-25 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1389 N$2778 N$2777 "Straight Waveguide" sch_x=-25 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1390 N$2780 N$2779 "Straight Waveguide" sch_x=-25 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1391 N$2782 N$2781 "Straight Waveguide" sch_x=-25 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1392 N$2784 N$2783 "Straight Waveguide" sch_x=-25 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1393 N$2786 N$2785 "Straight Waveguide" sch_x=-25 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1394 N$2788 N$2787 "Straight Waveguide" sch_x=-25 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1395 N$2790 N$2789 "Straight Waveguide" sch_x=-25 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1396 N$2792 N$2791 "Straight Waveguide" sch_x=-25 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1397 N$2794 N$2793 "Straight Waveguide" sch_x=-23 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1398 N$2796 N$2795 "Straight Waveguide" sch_x=-23 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1399 N$2798 N$2797 "Straight Waveguide" sch_x=-23 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1400 N$2800 N$2799 "Straight Waveguide" sch_x=-23 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1401 N$2802 N$2801 "Straight Waveguide" sch_x=-23 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1402 N$2804 N$2803 "Straight Waveguide" sch_x=-23 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1403 N$2806 N$2805 "Straight Waveguide" sch_x=-23 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1404 N$2808 N$2807 "Straight Waveguide" sch_x=-23 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1405 N$2810 N$2809 "Straight Waveguide" sch_x=-21 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1406 N$2812 N$2811 "Straight Waveguide" sch_x=-21 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1407 N$2814 N$2813 "Straight Waveguide" sch_x=-21 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1408 N$2816 N$2815 "Straight Waveguide" sch_x=-21 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1409 N$2818 N$2817 "Straight Waveguide" sch_x=-21 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1410 N$2820 N$2819 "Straight Waveguide" sch_x=-21 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1411 N$2822 N$2821 "Straight Waveguide" sch_x=-19 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1412 N$2824 N$2823 "Straight Waveguide" sch_x=-19 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1413 N$2826 N$2825 "Straight Waveguide" sch_x=-19 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1414 N$2828 N$2827 "Straight Waveguide" sch_x=-19 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1415 N$2830 N$2829 "Straight Waveguide" sch_x=-17 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1416 N$2832 N$2831 "Straight Waveguide" sch_x=-17 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1417 N$2833 N$2834 "Straight Waveguide" sch_x=-21 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1418 N$2835 N$2836 "Straight Waveguide" sch_x=-20 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1419 N$2837 N$2838 "Straight Waveguide" sch_x=-19 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1420 N$2839 N$2840 "Straight Waveguide" sch_x=-18 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1421 N$2841 N$2842 "Straight Waveguide" sch_x=-17 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1422 N$2843 N$2844 "Straight Waveguide" sch_x=-16 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1423 N$2845 N$2846 "Straight Waveguide" sch_x=-15 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1424 N$2847 N$2848 "Straight Waveguide" sch_x=-15 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1425 N$2849 N$2850 "Straight Waveguide" sch_x=-16 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1426 N$2851 N$2852 "Straight Waveguide" sch_x=-17 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1427 N$2853 N$2854 "Straight Waveguide" sch_x=-18 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1428 N$2855 N$2856 "Straight Waveguide" sch_x=-19 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1429 N$2857 N$2858 "Straight Waveguide" sch_x=-20 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1430 N$2859 N$2860 "Straight Waveguide" sch_x=-21 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1431 N$2861 N$2862 "Straight Waveguide" sch_x=-22 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1432 N$2863 N$2864 "Straight Waveguide" sch_x=-22 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1433 N$2865 N$2866 "Straight Waveguide" sch_x=29 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1434 N$2867 N$2868 "Straight Waveguide" sch_x=29 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1435 N$2869 N$2870 "Straight Waveguide" sch_x=29 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1436 N$2871 N$2872 "Straight Waveguide" sch_x=29 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1437 N$2873 N$2874 "Straight Waveguide" sch_x=29 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1438 N$2875 N$2876 "Straight Waveguide" sch_x=29 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1439 N$2877 N$2878 "Straight Waveguide" sch_x=29 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1440 N$2879 N$2880 "Straight Waveguide" sch_x=29 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1441 N$2881 N$2882 "Straight Waveguide" sch_x=29 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1442 N$2883 N$2884 "Straight Waveguide" sch_x=29 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1443 N$2885 N$2886 "Straight Waveguide" sch_x=29 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1444 N$2887 N$2888 "Straight Waveguide" sch_x=29 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1445 N$2889 N$2890 "Straight Waveguide" sch_x=29 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1446 N$2891 N$2892 "Straight Waveguide" sch_x=29 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1447 N$2893 N$2894 "Straight Waveguide" sch_x=27 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1448 N$2895 N$2896 "Straight Waveguide" sch_x=27 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1449 N$2897 N$2898 "Straight Waveguide" sch_x=27 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1450 N$2899 N$2900 "Straight Waveguide" sch_x=27 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1451 N$2901 N$2902 "Straight Waveguide" sch_x=27 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1452 N$2903 N$2904 "Straight Waveguide" sch_x=27 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1453 N$2905 N$2906 "Straight Waveguide" sch_x=27 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1454 N$2907 N$2908 "Straight Waveguide" sch_x=27 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1455 N$2909 N$2910 "Straight Waveguide" sch_x=27 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1456 N$2911 N$2912 "Straight Waveguide" sch_x=27 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1457 N$2913 N$2914 "Straight Waveguide" sch_x=27 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1458 N$2915 N$2916 "Straight Waveguide" sch_x=27 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1459 N$2917 N$2918 "Straight Waveguide" sch_x=25 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1460 N$2919 N$2920 "Straight Waveguide" sch_x=25 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1461 N$2921 N$2922 "Straight Waveguide" sch_x=25 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1462 N$2923 N$2924 "Straight Waveguide" sch_x=25 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1463 N$2925 N$2926 "Straight Waveguide" sch_x=25 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1464 N$2927 N$2928 "Straight Waveguide" sch_x=25 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1465 N$2929 N$2930 "Straight Waveguide" sch_x=25 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1466 N$2931 N$2932 "Straight Waveguide" sch_x=25 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1467 N$2933 N$2934 "Straight Waveguide" sch_x=25 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1468 N$2935 N$2936 "Straight Waveguide" sch_x=25 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1469 N$2937 N$2938 "Straight Waveguide" sch_x=23 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1470 N$2939 N$2940 "Straight Waveguide" sch_x=23 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1471 N$2941 N$2942 "Straight Waveguide" sch_x=23 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1472 N$2943 N$2944 "Straight Waveguide" sch_x=23 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1473 N$2945 N$2946 "Straight Waveguide" sch_x=23 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1474 N$2947 N$2948 "Straight Waveguide" sch_x=23 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1475 N$2949 N$2950 "Straight Waveguide" sch_x=23 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1476 N$2951 N$2952 "Straight Waveguide" sch_x=23 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1477 N$2953 N$2954 "Straight Waveguide" sch_x=21 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1478 N$2955 N$2956 "Straight Waveguide" sch_x=21 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1479 N$2957 N$2958 "Straight Waveguide" sch_x=21 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1480 N$2959 N$2960 "Straight Waveguide" sch_x=21 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1481 N$2961 N$2962 "Straight Waveguide" sch_x=21 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1482 N$2963 N$2964 "Straight Waveguide" sch_x=21 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1483 N$2965 N$2966 "Straight Waveguide" sch_x=19 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1484 N$2967 N$2968 "Straight Waveguide" sch_x=19 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1485 N$2969 N$2970 "Straight Waveguide" sch_x=19 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1486 N$2971 N$2972 "Straight Waveguide" sch_x=19 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1487 N$2973 N$2974 "Straight Waveguide" sch_x=17 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1488 N$2975 N$2976 "Straight Waveguide" sch_x=17 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1489 N$2978 N$2977 "Straight Waveguide" sch_x=21 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1490 N$2980 N$2979 "Straight Waveguide" sch_x=20 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1491 N$2982 N$2981 "Straight Waveguide" sch_x=19 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1492 N$2984 N$2983 "Straight Waveguide" sch_x=18 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1493 N$2986 N$2985 "Straight Waveguide" sch_x=17 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1494 N$2988 N$2987 "Straight Waveguide" sch_x=16 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1495 N$2990 N$2989 "Straight Waveguide" sch_x=15 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1496 N$2992 N$2991 "Straight Waveguide" sch_x=15 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1497 N$2994 N$2993 "Straight Waveguide" sch_x=16 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1498 N$2996 N$2995 "Straight Waveguide" sch_x=17 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1499 N$2998 N$2997 "Straight Waveguide" sch_x=18 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1500 N$3000 N$2999 "Straight Waveguide" sch_x=19 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1501 N$3002 N$3001 "Straight Waveguide" sch_x=20 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1502 N$3004 N$3003 "Straight Waveguide" sch_x=21 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1503 N$3006 N$3005 "Straight Waveguide" sch_x=22 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1504 N$3008 N$3007 "Straight Waveguide" sch_x=22 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1505 N$3009 N$3010 "Straight Waveguide" sch_x=-4 sch_y=15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1506 N$3011 N$3012 "Straight Waveguide" sch_x=-5 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1507 N$3013 N$3014 "Straight Waveguide" sch_x=-5 sch_y=13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1508 N$3015 N$3016 "Straight Waveguide" sch_x=-3 sch_y=14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1509 N$3017 N$3018 "Straight Waveguide" sch_x=-3 sch_y=13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1510 N$3019 N$3020 "Straight Waveguide" sch_x=-4 sch_y=12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1511 N$3021 N$3022 "Straight Waveguide" sch_x=0 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1512 N$3023 N$3024 "Straight Waveguide" sch_x=-1 sch_y=15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1513 N$3025 N$3026 "Straight Waveguide" sch_x=-1 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1514 N$3027 N$3028 "Straight Waveguide" sch_x=1 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1515 N$3029 N$3030 "Straight Waveguide" sch_x=1 sch_y=15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1516 N$3031 N$3032 "Straight Waveguide" sch_x=0 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1517 N$3033 N$3034 "Straight Waveguide" sch_x=0 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1518 N$3035 N$3036 "Straight Waveguide" sch_x=-1 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1519 N$3037 N$3038 "Straight Waveguide" sch_x=-1 sch_y=12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1520 N$3039 N$3040 "Straight Waveguide" sch_x=1 sch_y=12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1521 N$3041 N$3042 "Straight Waveguide" sch_x=1 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1522 N$3043 N$3044 "Straight Waveguide" sch_x=0 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1523 N$3045 N$3046 "Straight Waveguide" sch_x=4 sch_y=15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1524 N$3047 N$3048 "Straight Waveguide" sch_x=3 sch_y=14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1525 N$3049 N$3050 "Straight Waveguide" sch_x=3 sch_y=13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1526 N$3051 N$3052 "Straight Waveguide" sch_x=5 sch_y=13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1527 N$3053 N$3054 "Straight Waveguide" sch_x=5 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1528 N$3055 N$3056 "Straight Waveguide" sch_x=4 sch_y=12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1529 N$3057 N$3058 "Straight Waveguide" sch_x=-4 sch_y=11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1530 N$3059 N$3060 "Straight Waveguide" sch_x=-5 sch_y=10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1531 N$3061 N$3062 "Straight Waveguide" sch_x=-5 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1532 N$3063 N$3064 "Straight Waveguide" sch_x=-3 sch_y=10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1533 N$3065 N$3066 "Straight Waveguide" sch_x=-3 sch_y=9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1534 N$3067 N$3068 "Straight Waveguide" sch_x=-4 sch_y=8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1535 N$3069 N$3070 "Straight Waveguide" sch_x=0 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1536 N$3071 N$3072 "Straight Waveguide" sch_x=-1 sch_y=11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1537 N$3073 N$3074 "Straight Waveguide" sch_x=-1 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1538 N$3075 N$3076 "Straight Waveguide" sch_x=1 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1539 N$3077 N$3078 "Straight Waveguide" sch_x=1 sch_y=11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1540 N$3079 N$3080 "Straight Waveguide" sch_x=0 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1541 N$3081 N$3082 "Straight Waveguide" sch_x=0 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1542 N$3083 N$3084 "Straight Waveguide" sch_x=-1 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1543 N$3085 N$3086 "Straight Waveguide" sch_x=-1 sch_y=8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1544 N$3087 N$3088 "Straight Waveguide" sch_x=1 sch_y=8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1545 N$3089 N$3090 "Straight Waveguide" sch_x=1 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1546 N$3091 N$3092 "Straight Waveguide" sch_x=0 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1547 N$3093 N$3094 "Straight Waveguide" sch_x=4 sch_y=11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1548 N$3095 N$3096 "Straight Waveguide" sch_x=3 sch_y=10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1549 N$3097 N$3098 "Straight Waveguide" sch_x=3 sch_y=9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1550 N$3099 N$3100 "Straight Waveguide" sch_x=5 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1551 N$3101 N$3102 "Straight Waveguide" sch_x=5 sch_y=10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1552 N$3103 N$3104 "Straight Waveguide" sch_x=4 sch_y=8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1553 N$3106 N$3105 "Straight Waveguide" sch_x=-13 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1554 N$3108 N$3107 "Straight Waveguide" sch_x=-13 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1555 N$3110 N$3109 "Straight Waveguide" sch_x=-13 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1556 N$3112 N$3111 "Straight Waveguide" sch_x=-13 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1557 N$3114 N$3113 "Straight Waveguide" sch_x=-13 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1558 N$3116 N$3115 "Straight Waveguide" sch_x=-13 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1559 N$3118 N$3117 "Straight Waveguide" sch_x=-11 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1560 N$3120 N$3119 "Straight Waveguide" sch_x=-11 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1561 N$3122 N$3121 "Straight Waveguide" sch_x=-11 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1562 N$3124 N$3123 "Straight Waveguide" sch_x=-11 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1563 N$3126 N$3125 "Straight Waveguide" sch_x=-9 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1564 N$3128 N$3127 "Straight Waveguide" sch_x=-9 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1565 N$3129 N$3130 "Straight Waveguide" sch_x=-9 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1566 N$3131 N$3132 "Straight Waveguide" sch_x=-8 sch_y=13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1567 N$3133 N$3134 "Straight Waveguide" sch_x=-7 sch_y=12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1568 N$3135 N$3136 "Straight Waveguide" sch_x=-7 sch_y=11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1569 N$3137 N$3138 "Straight Waveguide" sch_x=-8 sch_y=10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1570 N$3139 N$3140 "Straight Waveguide" sch_x=-9 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1571 N$3141 N$3142 "Straight Waveguide" sch_x=-10 sch_y=14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1572 N$3143 N$3144 "Straight Waveguide" sch_x=-10 sch_y=9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1573 N$3145 N$3146 "Straight Waveguide" sch_x=13 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1574 N$3147 N$3148 "Straight Waveguide" sch_x=13 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1575 N$3149 N$3150 "Straight Waveguide" sch_x=13 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1576 N$3151 N$3152 "Straight Waveguide" sch_x=13 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1577 N$3153 N$3154 "Straight Waveguide" sch_x=13 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1578 N$3155 N$3156 "Straight Waveguide" sch_x=13 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1579 N$3157 N$3158 "Straight Waveguide" sch_x=11 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1580 N$3159 N$3160 "Straight Waveguide" sch_x=11 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1581 N$3161 N$3162 "Straight Waveguide" sch_x=11 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1582 N$3163 N$3164 "Straight Waveguide" sch_x=11 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1583 N$3165 N$3166 "Straight Waveguide" sch_x=9 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1584 N$3167 N$3168 "Straight Waveguide" sch_x=9 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1585 N$3170 N$3169 "Straight Waveguide" sch_x=9 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1586 N$3172 N$3171 "Straight Waveguide" sch_x=8 sch_y=13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1587 N$3174 N$3173 "Straight Waveguide" sch_x=7 sch_y=12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1588 N$3176 N$3175 "Straight Waveguide" sch_x=7 sch_y=11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1589 N$3178 N$3177 "Straight Waveguide" sch_x=8 sch_y=10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1590 N$3180 N$3179 "Straight Waveguide" sch_x=9 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1591 N$3182 N$3181 "Straight Waveguide" sch_x=10 sch_y=14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1592 N$3184 N$3183 "Straight Waveguide" sch_x=10 sch_y=9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1593 N$3185 N$3186 "Straight Waveguide" sch_x=-4 sch_y=7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1594 N$3187 N$3188 "Straight Waveguide" sch_x=-5 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1595 N$3189 N$3190 "Straight Waveguide" sch_x=-5 sch_y=5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1596 N$3191 N$3192 "Straight Waveguide" sch_x=-3 sch_y=6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1597 N$3193 N$3194 "Straight Waveguide" sch_x=-3 sch_y=5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1598 N$3195 N$3196 "Straight Waveguide" sch_x=-4 sch_y=4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1599 N$3197 N$3198 "Straight Waveguide" sch_x=0 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1600 N$3199 N$3200 "Straight Waveguide" sch_x=-1 sch_y=7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1601 N$3201 N$3202 "Straight Waveguide" sch_x=-1 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1602 N$3203 N$3204 "Straight Waveguide" sch_x=1 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1603 N$3205 N$3206 "Straight Waveguide" sch_x=1 sch_y=7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1604 N$3207 N$3208 "Straight Waveguide" sch_x=0 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1605 N$3209 N$3210 "Straight Waveguide" sch_x=0 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1606 N$3211 N$3212 "Straight Waveguide" sch_x=-1 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1607 N$3213 N$3214 "Straight Waveguide" sch_x=-1 sch_y=4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1608 N$3215 N$3216 "Straight Waveguide" sch_x=1 sch_y=4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1609 N$3217 N$3218 "Straight Waveguide" sch_x=1 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1610 N$3219 N$3220 "Straight Waveguide" sch_x=0 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1611 N$3221 N$3222 "Straight Waveguide" sch_x=4 sch_y=7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1612 N$3223 N$3224 "Straight Waveguide" sch_x=3 sch_y=6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1613 N$3225 N$3226 "Straight Waveguide" sch_x=3 sch_y=5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1614 N$3227 N$3228 "Straight Waveguide" sch_x=5 sch_y=5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1615 N$3229 N$3230 "Straight Waveguide" sch_x=5 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1616 N$3231 N$3232 "Straight Waveguide" sch_x=4 sch_y=4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1617 N$3233 N$3234 "Straight Waveguide" sch_x=-4 sch_y=3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1618 N$3235 N$3236 "Straight Waveguide" sch_x=-5 sch_y=2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1619 N$3237 N$3238 "Straight Waveguide" sch_x=-5 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1620 N$3239 N$3240 "Straight Waveguide" sch_x=-3 sch_y=2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1621 N$3241 N$3242 "Straight Waveguide" sch_x=-3 sch_y=1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1622 N$3243 N$3244 "Straight Waveguide" sch_x=-4 sch_y=0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1623 N$3245 N$3246 "Straight Waveguide" sch_x=0 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1624 N$3247 N$3248 "Straight Waveguide" sch_x=-1 sch_y=3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1625 N$3249 N$3250 "Straight Waveguide" sch_x=-1 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1626 N$3251 N$3252 "Straight Waveguide" sch_x=1 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1627 N$3253 N$3254 "Straight Waveguide" sch_x=1 sch_y=3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1628 N$3255 N$3256 "Straight Waveguide" sch_x=0 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1629 N$3257 N$3258 "Straight Waveguide" sch_x=0 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1630 N$3259 N$3260 "Straight Waveguide" sch_x=-1 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1631 N$3261 N$3262 "Straight Waveguide" sch_x=-1 sch_y=0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1632 N$3263 N$3264 "Straight Waveguide" sch_x=1 sch_y=0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1633 N$3265 N$3266 "Straight Waveguide" sch_x=1 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1634 N$3267 N$3268 "Straight Waveguide" sch_x=0 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1635 N$3269 N$3270 "Straight Waveguide" sch_x=4 sch_y=3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1636 N$3271 N$3272 "Straight Waveguide" sch_x=3 sch_y=2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1637 N$3273 N$3274 "Straight Waveguide" sch_x=3 sch_y=1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1638 N$3275 N$3276 "Straight Waveguide" sch_x=5 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1639 N$3277 N$3278 "Straight Waveguide" sch_x=5 sch_y=2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1640 N$3279 N$3280 "Straight Waveguide" sch_x=4 sch_y=0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1641 N$3282 N$3281 "Straight Waveguide" sch_x=-13 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1642 N$3284 N$3283 "Straight Waveguide" sch_x=-13 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1643 N$3286 N$3285 "Straight Waveguide" sch_x=-13 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1644 N$3288 N$3287 "Straight Waveguide" sch_x=-13 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1645 N$3290 N$3289 "Straight Waveguide" sch_x=-13 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1646 N$3292 N$3291 "Straight Waveguide" sch_x=-13 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1647 N$3294 N$3293 "Straight Waveguide" sch_x=-11 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1648 N$3296 N$3295 "Straight Waveguide" sch_x=-11 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1649 N$3298 N$3297 "Straight Waveguide" sch_x=-11 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1650 N$3300 N$3299 "Straight Waveguide" sch_x=-11 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1651 N$3302 N$3301 "Straight Waveguide" sch_x=-9 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1652 N$3304 N$3303 "Straight Waveguide" sch_x=-9 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1653 N$3305 N$3306 "Straight Waveguide" sch_x=-9 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1654 N$3307 N$3308 "Straight Waveguide" sch_x=-8 sch_y=5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1655 N$3309 N$3310 "Straight Waveguide" sch_x=-7 sch_y=4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1656 N$3311 N$3312 "Straight Waveguide" sch_x=-7 sch_y=3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1657 N$3313 N$3314 "Straight Waveguide" sch_x=-8 sch_y=2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1658 N$3315 N$3316 "Straight Waveguide" sch_x=-9 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1659 N$3317 N$3318 "Straight Waveguide" sch_x=-10 sch_y=6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1660 N$3319 N$3320 "Straight Waveguide" sch_x=-10 sch_y=1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1661 N$3321 N$3322 "Straight Waveguide" sch_x=13 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1662 N$3323 N$3324 "Straight Waveguide" sch_x=13 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1663 N$3325 N$3326 "Straight Waveguide" sch_x=13 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1664 N$3327 N$3328 "Straight Waveguide" sch_x=13 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1665 N$3329 N$3330 "Straight Waveguide" sch_x=13 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1666 N$3331 N$3332 "Straight Waveguide" sch_x=13 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1667 N$3333 N$3334 "Straight Waveguide" sch_x=11 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1668 N$3335 N$3336 "Straight Waveguide" sch_x=11 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1669 N$3337 N$3338 "Straight Waveguide" sch_x=11 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1670 N$3339 N$3340 "Straight Waveguide" sch_x=11 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1671 N$3341 N$3342 "Straight Waveguide" sch_x=9 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1672 N$3343 N$3344 "Straight Waveguide" sch_x=9 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1673 N$3346 N$3345 "Straight Waveguide" sch_x=9 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1674 N$3348 N$3347 "Straight Waveguide" sch_x=8 sch_y=5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1675 N$3350 N$3349 "Straight Waveguide" sch_x=7 sch_y=4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1676 N$3352 N$3351 "Straight Waveguide" sch_x=7 sch_y=3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1677 N$3354 N$3353 "Straight Waveguide" sch_x=8 sch_y=2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1678 N$3356 N$3355 "Straight Waveguide" sch_x=9 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1679 N$3358 N$3357 "Straight Waveguide" sch_x=10 sch_y=6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1680 N$3360 N$3359 "Straight Waveguide" sch_x=10 sch_y=1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1681 N$3362 N$3361 "Straight Waveguide" sch_x=-29 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1682 N$3364 N$3363 "Straight Waveguide" sch_x=-29 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1683 N$3366 N$3365 "Straight Waveguide" sch_x=-29 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1684 N$3368 N$3367 "Straight Waveguide" sch_x=-29 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1685 N$3370 N$3369 "Straight Waveguide" sch_x=-29 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1686 N$3372 N$3371 "Straight Waveguide" sch_x=-29 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1687 N$3374 N$3373 "Straight Waveguide" sch_x=-29 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1688 N$3376 N$3375 "Straight Waveguide" sch_x=-29 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1689 N$3378 N$3377 "Straight Waveguide" sch_x=-29 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1690 N$3380 N$3379 "Straight Waveguide" sch_x=-29 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1691 N$3382 N$3381 "Straight Waveguide" sch_x=-29 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1692 N$3384 N$3383 "Straight Waveguide" sch_x=-29 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1693 N$3386 N$3385 "Straight Waveguide" sch_x=-29 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1694 N$3388 N$3387 "Straight Waveguide" sch_x=-29 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1695 N$3390 N$3389 "Straight Waveguide" sch_x=-27 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1696 N$3392 N$3391 "Straight Waveguide" sch_x=-27 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1697 N$3394 N$3393 "Straight Waveguide" sch_x=-27 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1698 N$3396 N$3395 "Straight Waveguide" sch_x=-27 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1699 N$3398 N$3397 "Straight Waveguide" sch_x=-27 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1700 N$3400 N$3399 "Straight Waveguide" sch_x=-27 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1701 N$3402 N$3401 "Straight Waveguide" sch_x=-27 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1702 N$3404 N$3403 "Straight Waveguide" sch_x=-27 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1703 N$3406 N$3405 "Straight Waveguide" sch_x=-27 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1704 N$3408 N$3407 "Straight Waveguide" sch_x=-27 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1705 N$3410 N$3409 "Straight Waveguide" sch_x=-27 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1706 N$3412 N$3411 "Straight Waveguide" sch_x=-27 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1707 N$3414 N$3413 "Straight Waveguide" sch_x=-25 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1708 N$3416 N$3415 "Straight Waveguide" sch_x=-25 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1709 N$3418 N$3417 "Straight Waveguide" sch_x=-25 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1710 N$3420 N$3419 "Straight Waveguide" sch_x=-25 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1711 N$3422 N$3421 "Straight Waveguide" sch_x=-25 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1712 N$3424 N$3423 "Straight Waveguide" sch_x=-25 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1713 N$3426 N$3425 "Straight Waveguide" sch_x=-25 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1714 N$3428 N$3427 "Straight Waveguide" sch_x=-25 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1715 N$3430 N$3429 "Straight Waveguide" sch_x=-25 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1716 N$3432 N$3431 "Straight Waveguide" sch_x=-25 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1717 N$3434 N$3433 "Straight Waveguide" sch_x=-23 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1718 N$3436 N$3435 "Straight Waveguide" sch_x=-23 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1719 N$3438 N$3437 "Straight Waveguide" sch_x=-23 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1720 N$3440 N$3439 "Straight Waveguide" sch_x=-23 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1721 N$3442 N$3441 "Straight Waveguide" sch_x=-23 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1722 N$3444 N$3443 "Straight Waveguide" sch_x=-23 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1723 N$3446 N$3445 "Straight Waveguide" sch_x=-23 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1724 N$3448 N$3447 "Straight Waveguide" sch_x=-23 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1725 N$3450 N$3449 "Straight Waveguide" sch_x=-21 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1726 N$3452 N$3451 "Straight Waveguide" sch_x=-21 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1727 N$3454 N$3453 "Straight Waveguide" sch_x=-21 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1728 N$3456 N$3455 "Straight Waveguide" sch_x=-21 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1729 N$3458 N$3457 "Straight Waveguide" sch_x=-21 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1730 N$3460 N$3459 "Straight Waveguide" sch_x=-21 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1731 N$3462 N$3461 "Straight Waveguide" sch_x=-19 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1732 N$3464 N$3463 "Straight Waveguide" sch_x=-19 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1733 N$3466 N$3465 "Straight Waveguide" sch_x=-19 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1734 N$3468 N$3467 "Straight Waveguide" sch_x=-19 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1735 N$3470 N$3469 "Straight Waveguide" sch_x=-17 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1736 N$3472 N$3471 "Straight Waveguide" sch_x=-17 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1737 N$3473 N$3474 "Straight Waveguide" sch_x=-21 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1738 N$3475 N$3476 "Straight Waveguide" sch_x=-20 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1739 N$3477 N$3478 "Straight Waveguide" sch_x=-19 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1740 N$3479 N$3480 "Straight Waveguide" sch_x=-18 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1741 N$3481 N$3482 "Straight Waveguide" sch_x=-17 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1742 N$3483 N$3484 "Straight Waveguide" sch_x=-16 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1743 N$3485 N$3486 "Straight Waveguide" sch_x=-15 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1744 N$3487 N$3488 "Straight Waveguide" sch_x=-15 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1745 N$3489 N$3490 "Straight Waveguide" sch_x=-16 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1746 N$3491 N$3492 "Straight Waveguide" sch_x=-17 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1747 N$3493 N$3494 "Straight Waveguide" sch_x=-18 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1748 N$3495 N$3496 "Straight Waveguide" sch_x=-19 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1749 N$3497 N$3498 "Straight Waveguide" sch_x=-20 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1750 N$3499 N$3500 "Straight Waveguide" sch_x=-21 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1751 N$3501 N$3502 "Straight Waveguide" sch_x=-22 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1752 N$3503 N$3504 "Straight Waveguide" sch_x=-22 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1753 N$3505 N$3506 "Straight Waveguide" sch_x=29 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1754 N$3507 N$3508 "Straight Waveguide" sch_x=29 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1755 N$3509 N$3510 "Straight Waveguide" sch_x=29 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1756 N$3511 N$3512 "Straight Waveguide" sch_x=29 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1757 N$3513 N$3514 "Straight Waveguide" sch_x=29 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1758 N$3515 N$3516 "Straight Waveguide" sch_x=29 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1759 N$3517 N$3518 "Straight Waveguide" sch_x=29 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1760 N$3519 N$3520 "Straight Waveguide" sch_x=29 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1761 N$3521 N$3522 "Straight Waveguide" sch_x=29 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1762 N$3523 N$3524 "Straight Waveguide" sch_x=29 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1763 N$3525 N$3526 "Straight Waveguide" sch_x=29 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1764 N$3527 N$3528 "Straight Waveguide" sch_x=29 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1765 N$3529 N$3530 "Straight Waveguide" sch_x=29 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1766 N$3531 N$3532 "Straight Waveguide" sch_x=29 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1767 N$3533 N$3534 "Straight Waveguide" sch_x=27 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1768 N$3535 N$3536 "Straight Waveguide" sch_x=27 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1769 N$3537 N$3538 "Straight Waveguide" sch_x=27 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1770 N$3539 N$3540 "Straight Waveguide" sch_x=27 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1771 N$3541 N$3542 "Straight Waveguide" sch_x=27 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1772 N$3543 N$3544 "Straight Waveguide" sch_x=27 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1773 N$3545 N$3546 "Straight Waveguide" sch_x=27 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1774 N$3547 N$3548 "Straight Waveguide" sch_x=27 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1775 N$3549 N$3550 "Straight Waveguide" sch_x=27 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1776 N$3551 N$3552 "Straight Waveguide" sch_x=27 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1777 N$3553 N$3554 "Straight Waveguide" sch_x=27 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1778 N$3555 N$3556 "Straight Waveguide" sch_x=27 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1779 N$3557 N$3558 "Straight Waveguide" sch_x=25 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1780 N$3559 N$3560 "Straight Waveguide" sch_x=25 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1781 N$3561 N$3562 "Straight Waveguide" sch_x=25 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1782 N$3563 N$3564 "Straight Waveguide" sch_x=25 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1783 N$3565 N$3566 "Straight Waveguide" sch_x=25 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1784 N$3567 N$3568 "Straight Waveguide" sch_x=25 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1785 N$3569 N$3570 "Straight Waveguide" sch_x=25 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1786 N$3571 N$3572 "Straight Waveguide" sch_x=25 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1787 N$3573 N$3574 "Straight Waveguide" sch_x=25 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1788 N$3575 N$3576 "Straight Waveguide" sch_x=25 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1789 N$3577 N$3578 "Straight Waveguide" sch_x=23 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1790 N$3579 N$3580 "Straight Waveguide" sch_x=23 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1791 N$3581 N$3582 "Straight Waveguide" sch_x=23 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1792 N$3583 N$3584 "Straight Waveguide" sch_x=23 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1793 N$3585 N$3586 "Straight Waveguide" sch_x=23 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1794 N$3587 N$3588 "Straight Waveguide" sch_x=23 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1795 N$3589 N$3590 "Straight Waveguide" sch_x=23 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1796 N$3591 N$3592 "Straight Waveguide" sch_x=23 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1797 N$3593 N$3594 "Straight Waveguide" sch_x=21 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1798 N$3595 N$3596 "Straight Waveguide" sch_x=21 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1799 N$3597 N$3598 "Straight Waveguide" sch_x=21 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1800 N$3599 N$3600 "Straight Waveguide" sch_x=21 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1801 N$3601 N$3602 "Straight Waveguide" sch_x=21 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1802 N$3603 N$3604 "Straight Waveguide" sch_x=21 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1803 N$3605 N$3606 "Straight Waveguide" sch_x=19 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1804 N$3607 N$3608 "Straight Waveguide" sch_x=19 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1805 N$3609 N$3610 "Straight Waveguide" sch_x=19 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1806 N$3611 N$3612 "Straight Waveguide" sch_x=19 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1807 N$3613 N$3614 "Straight Waveguide" sch_x=17 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1808 N$3615 N$3616 "Straight Waveguide" sch_x=17 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1809 N$3618 N$3617 "Straight Waveguide" sch_x=21 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1810 N$3620 N$3619 "Straight Waveguide" sch_x=20 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1811 N$3622 N$3621 "Straight Waveguide" sch_x=19 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1812 N$3624 N$3623 "Straight Waveguide" sch_x=18 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1813 N$3626 N$3625 "Straight Waveguide" sch_x=17 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1814 N$3628 N$3627 "Straight Waveguide" sch_x=16 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1815 N$3630 N$3629 "Straight Waveguide" sch_x=15 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1816 N$3632 N$3631 "Straight Waveguide" sch_x=15 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1817 N$3634 N$3633 "Straight Waveguide" sch_x=16 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1818 N$3636 N$3635 "Straight Waveguide" sch_x=17 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1819 N$3638 N$3637 "Straight Waveguide" sch_x=18 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1820 N$3640 N$3639 "Straight Waveguide" sch_x=19 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1821 N$3642 N$3641 "Straight Waveguide" sch_x=20 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1822 N$3644 N$3643 "Straight Waveguide" sch_x=21 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1823 N$3646 N$3645 "Straight Waveguide" sch_x=22 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1824 N$3648 N$3647 "Straight Waveguide" sch_x=22 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1825 N$3650 N$3649 "Straight Waveguide" sch_x=-61 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1826 N$3652 N$3651 "Straight Waveguide" sch_x=-61 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1827 N$3654 N$3653 "Straight Waveguide" sch_x=-61 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1828 N$3656 N$3655 "Straight Waveguide" sch_x=-61 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1829 N$3658 N$3657 "Straight Waveguide" sch_x=-61 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1830 N$3660 N$3659 "Straight Waveguide" sch_x=-61 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1831 N$3662 N$3661 "Straight Waveguide" sch_x=-61 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1832 N$3664 N$3663 "Straight Waveguide" sch_x=-61 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1833 N$3666 N$3665 "Straight Waveguide" sch_x=-61 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1834 N$3668 N$3667 "Straight Waveguide" sch_x=-61 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1835 N$3670 N$3669 "Straight Waveguide" sch_x=-61 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1836 N$3672 N$3671 "Straight Waveguide" sch_x=-61 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1837 N$3674 N$3673 "Straight Waveguide" sch_x=-61 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1838 N$3676 N$3675 "Straight Waveguide" sch_x=-61 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1839 N$3678 N$3677 "Straight Waveguide" sch_x=-61 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1840 N$3680 N$3679 "Straight Waveguide" sch_x=-61 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1841 N$3682 N$3681 "Straight Waveguide" sch_x=-61 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1842 N$3684 N$3683 "Straight Waveguide" sch_x=-61 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1843 N$3686 N$3685 "Straight Waveguide" sch_x=-61 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1844 N$3688 N$3687 "Straight Waveguide" sch_x=-61 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1845 N$3690 N$3689 "Straight Waveguide" sch_x=-61 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1846 N$3692 N$3691 "Straight Waveguide" sch_x=-61 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1847 N$3694 N$3693 "Straight Waveguide" sch_x=-61 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1848 N$3696 N$3695 "Straight Waveguide" sch_x=-61 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1849 N$3698 N$3697 "Straight Waveguide" sch_x=-61 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1850 N$3700 N$3699 "Straight Waveguide" sch_x=-61 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1851 N$3702 N$3701 "Straight Waveguide" sch_x=-61 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1852 N$3704 N$3703 "Straight Waveguide" sch_x=-61 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1853 N$3706 N$3705 "Straight Waveguide" sch_x=-61 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1854 N$3708 N$3707 "Straight Waveguide" sch_x=-61 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1855 N$3710 N$3709 "Straight Waveguide" sch_x=-59 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1856 N$3712 N$3711 "Straight Waveguide" sch_x=-59 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1857 N$3714 N$3713 "Straight Waveguide" sch_x=-59 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1858 N$3716 N$3715 "Straight Waveguide" sch_x=-59 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1859 N$3718 N$3717 "Straight Waveguide" sch_x=-59 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1860 N$3720 N$3719 "Straight Waveguide" sch_x=-59 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1861 N$3722 N$3721 "Straight Waveguide" sch_x=-59 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1862 N$3724 N$3723 "Straight Waveguide" sch_x=-59 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1863 N$3726 N$3725 "Straight Waveguide" sch_x=-59 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1864 N$3728 N$3727 "Straight Waveguide" sch_x=-59 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1865 N$3730 N$3729 "Straight Waveguide" sch_x=-59 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1866 N$3732 N$3731 "Straight Waveguide" sch_x=-59 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1867 N$3734 N$3733 "Straight Waveguide" sch_x=-59 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1868 N$3736 N$3735 "Straight Waveguide" sch_x=-59 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1869 N$3738 N$3737 "Straight Waveguide" sch_x=-59 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1870 N$3740 N$3739 "Straight Waveguide" sch_x=-59 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1871 N$3742 N$3741 "Straight Waveguide" sch_x=-59 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1872 N$3744 N$3743 "Straight Waveguide" sch_x=-59 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1873 N$3746 N$3745 "Straight Waveguide" sch_x=-59 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1874 N$3748 N$3747 "Straight Waveguide" sch_x=-59 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1875 N$3750 N$3749 "Straight Waveguide" sch_x=-59 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1876 N$3752 N$3751 "Straight Waveguide" sch_x=-59 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1877 N$3754 N$3753 "Straight Waveguide" sch_x=-59 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1878 N$3756 N$3755 "Straight Waveguide" sch_x=-59 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1879 N$3758 N$3757 "Straight Waveguide" sch_x=-59 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1880 N$3760 N$3759 "Straight Waveguide" sch_x=-59 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1881 N$3762 N$3761 "Straight Waveguide" sch_x=-59 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1882 N$3764 N$3763 "Straight Waveguide" sch_x=-59 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1883 N$3766 N$3765 "Straight Waveguide" sch_x=-57 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1884 N$3768 N$3767 "Straight Waveguide" sch_x=-57 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1885 N$3770 N$3769 "Straight Waveguide" sch_x=-57 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1886 N$3772 N$3771 "Straight Waveguide" sch_x=-57 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1887 N$3774 N$3773 "Straight Waveguide" sch_x=-57 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1888 N$3776 N$3775 "Straight Waveguide" sch_x=-57 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1889 N$3778 N$3777 "Straight Waveguide" sch_x=-57 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1890 N$3780 N$3779 "Straight Waveguide" sch_x=-57 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1891 N$3782 N$3781 "Straight Waveguide" sch_x=-57 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1892 N$3784 N$3783 "Straight Waveguide" sch_x=-57 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1893 N$3786 N$3785 "Straight Waveguide" sch_x=-57 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1894 N$3788 N$3787 "Straight Waveguide" sch_x=-57 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1895 N$3790 N$3789 "Straight Waveguide" sch_x=-57 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1896 N$3792 N$3791 "Straight Waveguide" sch_x=-57 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1897 N$3794 N$3793 "Straight Waveguide" sch_x=-57 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1898 N$3796 N$3795 "Straight Waveguide" sch_x=-57 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1899 N$3798 N$3797 "Straight Waveguide" sch_x=-57 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1900 N$3800 N$3799 "Straight Waveguide" sch_x=-57 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1901 N$3802 N$3801 "Straight Waveguide" sch_x=-57 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1902 N$3804 N$3803 "Straight Waveguide" sch_x=-57 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1903 N$3806 N$3805 "Straight Waveguide" sch_x=-57 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1904 N$3808 N$3807 "Straight Waveguide" sch_x=-57 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1905 N$3810 N$3809 "Straight Waveguide" sch_x=-57 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1906 N$3812 N$3811 "Straight Waveguide" sch_x=-57 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1907 N$3814 N$3813 "Straight Waveguide" sch_x=-57 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1908 N$3816 N$3815 "Straight Waveguide" sch_x=-57 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1909 N$3818 N$3817 "Straight Waveguide" sch_x=-55 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1910 N$3820 N$3819 "Straight Waveguide" sch_x=-55 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1911 N$3822 N$3821 "Straight Waveguide" sch_x=-55 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1912 N$3824 N$3823 "Straight Waveguide" sch_x=-55 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1913 N$3826 N$3825 "Straight Waveguide" sch_x=-55 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1914 N$3828 N$3827 "Straight Waveguide" sch_x=-55 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1915 N$3830 N$3829 "Straight Waveguide" sch_x=-55 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1916 N$3832 N$3831 "Straight Waveguide" sch_x=-55 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1917 N$3834 N$3833 "Straight Waveguide" sch_x=-55 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1918 N$3836 N$3835 "Straight Waveguide" sch_x=-55 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1919 N$3838 N$3837 "Straight Waveguide" sch_x=-55 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1920 N$3840 N$3839 "Straight Waveguide" sch_x=-55 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1921 N$3842 N$3841 "Straight Waveguide" sch_x=-55 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1922 N$3844 N$3843 "Straight Waveguide" sch_x=-55 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1923 N$3846 N$3845 "Straight Waveguide" sch_x=-55 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1924 N$3848 N$3847 "Straight Waveguide" sch_x=-55 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1925 N$3850 N$3849 "Straight Waveguide" sch_x=-55 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1926 N$3852 N$3851 "Straight Waveguide" sch_x=-55 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1927 N$3854 N$3853 "Straight Waveguide" sch_x=-55 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1928 N$3856 N$3855 "Straight Waveguide" sch_x=-55 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1929 N$3858 N$3857 "Straight Waveguide" sch_x=-55 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1930 N$3860 N$3859 "Straight Waveguide" sch_x=-55 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1931 N$3862 N$3861 "Straight Waveguide" sch_x=-55 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1932 N$3864 N$3863 "Straight Waveguide" sch_x=-55 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1933 N$3866 N$3865 "Straight Waveguide" sch_x=-53 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1934 N$3868 N$3867 "Straight Waveguide" sch_x=-53 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1935 N$3870 N$3869 "Straight Waveguide" sch_x=-53 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1936 N$3872 N$3871 "Straight Waveguide" sch_x=-53 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1937 N$3874 N$3873 "Straight Waveguide" sch_x=-53 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1938 N$3876 N$3875 "Straight Waveguide" sch_x=-53 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1939 N$3878 N$3877 "Straight Waveguide" sch_x=-53 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1940 N$3880 N$3879 "Straight Waveguide" sch_x=-53 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1941 N$3882 N$3881 "Straight Waveguide" sch_x=-53 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1942 N$3884 N$3883 "Straight Waveguide" sch_x=-53 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1943 N$3886 N$3885 "Straight Waveguide" sch_x=-53 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1944 N$3888 N$3887 "Straight Waveguide" sch_x=-53 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1945 N$3890 N$3889 "Straight Waveguide" sch_x=-53 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1946 N$3892 N$3891 "Straight Waveguide" sch_x=-53 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1947 N$3894 N$3893 "Straight Waveguide" sch_x=-53 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1948 N$3896 N$3895 "Straight Waveguide" sch_x=-53 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1949 N$3898 N$3897 "Straight Waveguide" sch_x=-53 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1950 N$3900 N$3899 "Straight Waveguide" sch_x=-53 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1951 N$3902 N$3901 "Straight Waveguide" sch_x=-53 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1952 N$3904 N$3903 "Straight Waveguide" sch_x=-53 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1953 N$3906 N$3905 "Straight Waveguide" sch_x=-53 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1954 N$3908 N$3907 "Straight Waveguide" sch_x=-53 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1955 N$3910 N$3909 "Straight Waveguide" sch_x=-51 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1956 N$3912 N$3911 "Straight Waveguide" sch_x=-51 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1957 N$3914 N$3913 "Straight Waveguide" sch_x=-51 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1958 N$3916 N$3915 "Straight Waveguide" sch_x=-51 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1959 N$3918 N$3917 "Straight Waveguide" sch_x=-51 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1960 N$3920 N$3919 "Straight Waveguide" sch_x=-51 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1961 N$3922 N$3921 "Straight Waveguide" sch_x=-51 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1962 N$3924 N$3923 "Straight Waveguide" sch_x=-51 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1963 N$3926 N$3925 "Straight Waveguide" sch_x=-51 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1964 N$3928 N$3927 "Straight Waveguide" sch_x=-51 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1965 N$3930 N$3929 "Straight Waveguide" sch_x=-51 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1966 N$3932 N$3931 "Straight Waveguide" sch_x=-51 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1967 N$3934 N$3933 "Straight Waveguide" sch_x=-51 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1968 N$3936 N$3935 "Straight Waveguide" sch_x=-51 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1969 N$3938 N$3937 "Straight Waveguide" sch_x=-51 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1970 N$3940 N$3939 "Straight Waveguide" sch_x=-51 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1971 N$3942 N$3941 "Straight Waveguide" sch_x=-51 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1972 N$3944 N$3943 "Straight Waveguide" sch_x=-51 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1973 N$3946 N$3945 "Straight Waveguide" sch_x=-51 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1974 N$3948 N$3947 "Straight Waveguide" sch_x=-51 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1975 N$3950 N$3949 "Straight Waveguide" sch_x=-49 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1976 N$3952 N$3951 "Straight Waveguide" sch_x=-49 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1977 N$3954 N$3953 "Straight Waveguide" sch_x=-49 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1978 N$3956 N$3955 "Straight Waveguide" sch_x=-49 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1979 N$3958 N$3957 "Straight Waveguide" sch_x=-49 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1980 N$3960 N$3959 "Straight Waveguide" sch_x=-49 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1981 N$3962 N$3961 "Straight Waveguide" sch_x=-49 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1982 N$3964 N$3963 "Straight Waveguide" sch_x=-49 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1983 N$3966 N$3965 "Straight Waveguide" sch_x=-49 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1984 N$3968 N$3967 "Straight Waveguide" sch_x=-49 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1985 N$3970 N$3969 "Straight Waveguide" sch_x=-49 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1986 N$3972 N$3971 "Straight Waveguide" sch_x=-49 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1987 N$3974 N$3973 "Straight Waveguide" sch_x=-49 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1988 N$3976 N$3975 "Straight Waveguide" sch_x=-49 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1989 N$3978 N$3977 "Straight Waveguide" sch_x=-49 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1990 N$3980 N$3979 "Straight Waveguide" sch_x=-49 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1991 N$3982 N$3981 "Straight Waveguide" sch_x=-49 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1992 N$3984 N$3983 "Straight Waveguide" sch_x=-49 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1993 N$3986 N$3985 "Straight Waveguide" sch_x=-47 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1994 N$3988 N$3987 "Straight Waveguide" sch_x=-47 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1995 N$3990 N$3989 "Straight Waveguide" sch_x=-47 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1996 N$3992 N$3991 "Straight Waveguide" sch_x=-47 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1997 N$3994 N$3993 "Straight Waveguide" sch_x=-47 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1998 N$3996 N$3995 "Straight Waveguide" sch_x=-47 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1999 N$3998 N$3997 "Straight Waveguide" sch_x=-47 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2000 N$4000 N$3999 "Straight Waveguide" sch_x=-47 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2001 N$4002 N$4001 "Straight Waveguide" sch_x=-47 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2002 N$4004 N$4003 "Straight Waveguide" sch_x=-47 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2003 N$4006 N$4005 "Straight Waveguide" sch_x=-47 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2004 N$4008 N$4007 "Straight Waveguide" sch_x=-47 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2005 N$4010 N$4009 "Straight Waveguide" sch_x=-47 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2006 N$4012 N$4011 "Straight Waveguide" sch_x=-47 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2007 N$4014 N$4013 "Straight Waveguide" sch_x=-47 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2008 N$4016 N$4015 "Straight Waveguide" sch_x=-47 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2009 N$4018 N$4017 "Straight Waveguide" sch_x=-45 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2010 N$4020 N$4019 "Straight Waveguide" sch_x=-45 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2011 N$4022 N$4021 "Straight Waveguide" sch_x=-45 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2012 N$4024 N$4023 "Straight Waveguide" sch_x=-45 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2013 N$4026 N$4025 "Straight Waveguide" sch_x=-45 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2014 N$4028 N$4027 "Straight Waveguide" sch_x=-45 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2015 N$4030 N$4029 "Straight Waveguide" sch_x=-45 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2016 N$4032 N$4031 "Straight Waveguide" sch_x=-45 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2017 N$4034 N$4033 "Straight Waveguide" sch_x=-45 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2018 N$4036 N$4035 "Straight Waveguide" sch_x=-45 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2019 N$4038 N$4037 "Straight Waveguide" sch_x=-45 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2020 N$4040 N$4039 "Straight Waveguide" sch_x=-45 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2021 N$4042 N$4041 "Straight Waveguide" sch_x=-45 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2022 N$4044 N$4043 "Straight Waveguide" sch_x=-45 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2023 N$4046 N$4045 "Straight Waveguide" sch_x=-43 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2024 N$4048 N$4047 "Straight Waveguide" sch_x=-43 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2025 N$4050 N$4049 "Straight Waveguide" sch_x=-43 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2026 N$4052 N$4051 "Straight Waveguide" sch_x=-43 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2027 N$4054 N$4053 "Straight Waveguide" sch_x=-43 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2028 N$4056 N$4055 "Straight Waveguide" sch_x=-43 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2029 N$4058 N$4057 "Straight Waveguide" sch_x=-43 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2030 N$4060 N$4059 "Straight Waveguide" sch_x=-43 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2031 N$4062 N$4061 "Straight Waveguide" sch_x=-43 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2032 N$4064 N$4063 "Straight Waveguide" sch_x=-43 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2033 N$4066 N$4065 "Straight Waveguide" sch_x=-43 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2034 N$4068 N$4067 "Straight Waveguide" sch_x=-43 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2035 N$4070 N$4069 "Straight Waveguide" sch_x=-41 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2036 N$4072 N$4071 "Straight Waveguide" sch_x=-41 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2037 N$4074 N$4073 "Straight Waveguide" sch_x=-41 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2038 N$4076 N$4075 "Straight Waveguide" sch_x=-41 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2039 N$4078 N$4077 "Straight Waveguide" sch_x=-41 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2040 N$4080 N$4079 "Straight Waveguide" sch_x=-41 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2041 N$4082 N$4081 "Straight Waveguide" sch_x=-41 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2042 N$4084 N$4083 "Straight Waveguide" sch_x=-41 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2043 N$4086 N$4085 "Straight Waveguide" sch_x=-41 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2044 N$4088 N$4087 "Straight Waveguide" sch_x=-41 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2045 N$4090 N$4089 "Straight Waveguide" sch_x=-39 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2046 N$4092 N$4091 "Straight Waveguide" sch_x=-39 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2047 N$4094 N$4093 "Straight Waveguide" sch_x=-39 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2048 N$4096 N$4095 "Straight Waveguide" sch_x=-39 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2049 N$4098 N$4097 "Straight Waveguide" sch_x=-39 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2050 N$4100 N$4099 "Straight Waveguide" sch_x=-39 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2051 N$4102 N$4101 "Straight Waveguide" sch_x=-39 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2052 N$4104 N$4103 "Straight Waveguide" sch_x=-39 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2053 N$4106 N$4105 "Straight Waveguide" sch_x=-37 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2054 N$4108 N$4107 "Straight Waveguide" sch_x=-37 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2055 N$4110 N$4109 "Straight Waveguide" sch_x=-37 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2056 N$4112 N$4111 "Straight Waveguide" sch_x=-37 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2057 N$4114 N$4113 "Straight Waveguide" sch_x=-37 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2058 N$4116 N$4115 "Straight Waveguide" sch_x=-37 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2059 N$4118 N$4117 "Straight Waveguide" sch_x=-35 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2060 N$4120 N$4119 "Straight Waveguide" sch_x=-35 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2061 N$4122 N$4121 "Straight Waveguide" sch_x=-35 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2062 N$4124 N$4123 "Straight Waveguide" sch_x=-35 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2063 N$4126 N$4125 "Straight Waveguide" sch_x=-33 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2064 N$4128 N$4127 "Straight Waveguide" sch_x=-33 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2065 N$4129 N$4130 "Straight Waveguide" sch_x=-45 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2066 N$4131 N$4132 "Straight Waveguide" sch_x=-44 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2067 N$4133 N$4134 "Straight Waveguide" sch_x=-43 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2068 N$4135 N$4136 "Straight Waveguide" sch_x=-42 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2069 N$4137 N$4138 "Straight Waveguide" sch_x=-41 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2070 N$4139 N$4140 "Straight Waveguide" sch_x=-40 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2071 N$4141 N$4142 "Straight Waveguide" sch_x=-39 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2072 N$4143 N$4144 "Straight Waveguide" sch_x=-38 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2073 N$4145 N$4146 "Straight Waveguide" sch_x=-37 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2074 N$4147 N$4148 "Straight Waveguide" sch_x=-36 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2075 N$4149 N$4150 "Straight Waveguide" sch_x=-35 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2076 N$4151 N$4152 "Straight Waveguide" sch_x=-34 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2077 N$4153 N$4154 "Straight Waveguide" sch_x=-33 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2078 N$4155 N$4156 "Straight Waveguide" sch_x=-32 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2079 N$4157 N$4158 "Straight Waveguide" sch_x=-31 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2080 N$4159 N$4160 "Straight Waveguide" sch_x=-31 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2081 N$4161 N$4162 "Straight Waveguide" sch_x=-32 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2082 N$4163 N$4164 "Straight Waveguide" sch_x=-33 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2083 N$4165 N$4166 "Straight Waveguide" sch_x=-34 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2084 N$4167 N$4168 "Straight Waveguide" sch_x=-35 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2085 N$4169 N$4170 "Straight Waveguide" sch_x=-36 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2086 N$4171 N$4172 "Straight Waveguide" sch_x=-37 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2087 N$4173 N$4174 "Straight Waveguide" sch_x=-38 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2088 N$4175 N$4176 "Straight Waveguide" sch_x=-39 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2089 N$4177 N$4178 "Straight Waveguide" sch_x=-40 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2090 N$4179 N$4180 "Straight Waveguide" sch_x=-41 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2091 N$4181 N$4182 "Straight Waveguide" sch_x=-42 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2092 N$4183 N$4184 "Straight Waveguide" sch_x=-43 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2093 N$4185 N$4186 "Straight Waveguide" sch_x=-44 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2094 N$4187 N$4188 "Straight Waveguide" sch_x=-45 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2095 N$4189 N$4190 "Straight Waveguide" sch_x=-46 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2096 N$4191 N$4192 "Straight Waveguide" sch_x=-46 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2097 N$4193 N$4194 "Straight Waveguide" sch_x=61 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2098 N$4195 N$4196 "Straight Waveguide" sch_x=61 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2099 N$4197 N$4198 "Straight Waveguide" sch_x=61 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2100 N$4199 N$4200 "Straight Waveguide" sch_x=61 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2101 N$4201 N$4202 "Straight Waveguide" sch_x=61 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2102 N$4203 N$4204 "Straight Waveguide" sch_x=61 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2103 N$4205 N$4206 "Straight Waveguide" sch_x=61 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2104 N$4207 N$4208 "Straight Waveguide" sch_x=61 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2105 N$4209 N$4210 "Straight Waveguide" sch_x=61 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2106 N$4211 N$4212 "Straight Waveguide" sch_x=61 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2107 N$4213 N$4214 "Straight Waveguide" sch_x=61 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2108 N$4215 N$4216 "Straight Waveguide" sch_x=61 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2109 N$4217 N$4218 "Straight Waveguide" sch_x=61 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2110 N$4219 N$4220 "Straight Waveguide" sch_x=61 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2111 N$4221 N$4222 "Straight Waveguide" sch_x=61 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2112 N$4223 N$4224 "Straight Waveguide" sch_x=61 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2113 N$4225 N$4226 "Straight Waveguide" sch_x=61 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2114 N$4227 N$4228 "Straight Waveguide" sch_x=61 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2115 N$4229 N$4230 "Straight Waveguide" sch_x=61 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2116 N$4231 N$4232 "Straight Waveguide" sch_x=61 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2117 N$4233 N$4234 "Straight Waveguide" sch_x=61 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2118 N$4235 N$4236 "Straight Waveguide" sch_x=61 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2119 N$4237 N$4238 "Straight Waveguide" sch_x=61 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2120 N$4239 N$4240 "Straight Waveguide" sch_x=61 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2121 N$4241 N$4242 "Straight Waveguide" sch_x=61 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2122 N$4243 N$4244 "Straight Waveguide" sch_x=61 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2123 N$4245 N$4246 "Straight Waveguide" sch_x=61 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2124 N$4247 N$4248 "Straight Waveguide" sch_x=61 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2125 N$4249 N$4250 "Straight Waveguide" sch_x=61 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2126 N$4251 N$4252 "Straight Waveguide" sch_x=61 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2127 N$4253 N$4254 "Straight Waveguide" sch_x=59 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2128 N$4255 N$4256 "Straight Waveguide" sch_x=59 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2129 N$4257 N$4258 "Straight Waveguide" sch_x=59 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2130 N$4259 N$4260 "Straight Waveguide" sch_x=59 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2131 N$4261 N$4262 "Straight Waveguide" sch_x=59 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2132 N$4263 N$4264 "Straight Waveguide" sch_x=59 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2133 N$4265 N$4266 "Straight Waveguide" sch_x=59 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2134 N$4267 N$4268 "Straight Waveguide" sch_x=59 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2135 N$4269 N$4270 "Straight Waveguide" sch_x=59 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2136 N$4271 N$4272 "Straight Waveguide" sch_x=59 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2137 N$4273 N$4274 "Straight Waveguide" sch_x=59 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2138 N$4275 N$4276 "Straight Waveguide" sch_x=59 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2139 N$4277 N$4278 "Straight Waveguide" sch_x=59 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2140 N$4279 N$4280 "Straight Waveguide" sch_x=59 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2141 N$4281 N$4282 "Straight Waveguide" sch_x=59 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2142 N$4283 N$4284 "Straight Waveguide" sch_x=59 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2143 N$4285 N$4286 "Straight Waveguide" sch_x=59 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2144 N$4287 N$4288 "Straight Waveguide" sch_x=59 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2145 N$4289 N$4290 "Straight Waveguide" sch_x=59 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2146 N$4291 N$4292 "Straight Waveguide" sch_x=59 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2147 N$4293 N$4294 "Straight Waveguide" sch_x=59 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2148 N$4295 N$4296 "Straight Waveguide" sch_x=59 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2149 N$4297 N$4298 "Straight Waveguide" sch_x=59 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2150 N$4299 N$4300 "Straight Waveguide" sch_x=59 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2151 N$4301 N$4302 "Straight Waveguide" sch_x=59 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2152 N$4303 N$4304 "Straight Waveguide" sch_x=59 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2153 N$4305 N$4306 "Straight Waveguide" sch_x=59 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2154 N$4307 N$4308 "Straight Waveguide" sch_x=59 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2155 N$4309 N$4310 "Straight Waveguide" sch_x=57 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2156 N$4311 N$4312 "Straight Waveguide" sch_x=57 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2157 N$4313 N$4314 "Straight Waveguide" sch_x=57 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2158 N$4315 N$4316 "Straight Waveguide" sch_x=57 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2159 N$4317 N$4318 "Straight Waveguide" sch_x=57 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2160 N$4319 N$4320 "Straight Waveguide" sch_x=57 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2161 N$4321 N$4322 "Straight Waveguide" sch_x=57 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2162 N$4323 N$4324 "Straight Waveguide" sch_x=57 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2163 N$4325 N$4326 "Straight Waveguide" sch_x=57 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2164 N$4327 N$4328 "Straight Waveguide" sch_x=57 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2165 N$4329 N$4330 "Straight Waveguide" sch_x=57 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2166 N$4331 N$4332 "Straight Waveguide" sch_x=57 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2167 N$4333 N$4334 "Straight Waveguide" sch_x=57 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2168 N$4335 N$4336 "Straight Waveguide" sch_x=57 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2169 N$4337 N$4338 "Straight Waveguide" sch_x=57 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2170 N$4339 N$4340 "Straight Waveguide" sch_x=57 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2171 N$4341 N$4342 "Straight Waveguide" sch_x=57 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2172 N$4343 N$4344 "Straight Waveguide" sch_x=57 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2173 N$4345 N$4346 "Straight Waveguide" sch_x=57 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2174 N$4347 N$4348 "Straight Waveguide" sch_x=57 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2175 N$4349 N$4350 "Straight Waveguide" sch_x=57 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2176 N$4351 N$4352 "Straight Waveguide" sch_x=57 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2177 N$4353 N$4354 "Straight Waveguide" sch_x=57 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2178 N$4355 N$4356 "Straight Waveguide" sch_x=57 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2179 N$4357 N$4358 "Straight Waveguide" sch_x=57 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2180 N$4359 N$4360 "Straight Waveguide" sch_x=57 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2181 N$4361 N$4362 "Straight Waveguide" sch_x=55 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2182 N$4363 N$4364 "Straight Waveguide" sch_x=55 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2183 N$4365 N$4366 "Straight Waveguide" sch_x=55 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2184 N$4367 N$4368 "Straight Waveguide" sch_x=55 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2185 N$4369 N$4370 "Straight Waveguide" sch_x=55 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2186 N$4371 N$4372 "Straight Waveguide" sch_x=55 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2187 N$4373 N$4374 "Straight Waveguide" sch_x=55 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2188 N$4375 N$4376 "Straight Waveguide" sch_x=55 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2189 N$4377 N$4378 "Straight Waveguide" sch_x=55 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2190 N$4379 N$4380 "Straight Waveguide" sch_x=55 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2191 N$4381 N$4382 "Straight Waveguide" sch_x=55 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2192 N$4383 N$4384 "Straight Waveguide" sch_x=55 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2193 N$4385 N$4386 "Straight Waveguide" sch_x=55 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2194 N$4387 N$4388 "Straight Waveguide" sch_x=55 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2195 N$4389 N$4390 "Straight Waveguide" sch_x=55 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2196 N$4391 N$4392 "Straight Waveguide" sch_x=55 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2197 N$4393 N$4394 "Straight Waveguide" sch_x=55 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2198 N$4395 N$4396 "Straight Waveguide" sch_x=55 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2199 N$4397 N$4398 "Straight Waveguide" sch_x=55 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2200 N$4399 N$4400 "Straight Waveguide" sch_x=55 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2201 N$4401 N$4402 "Straight Waveguide" sch_x=55 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2202 N$4403 N$4404 "Straight Waveguide" sch_x=55 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2203 N$4405 N$4406 "Straight Waveguide" sch_x=55 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2204 N$4407 N$4408 "Straight Waveguide" sch_x=55 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2205 N$4409 N$4410 "Straight Waveguide" sch_x=53 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2206 N$4411 N$4412 "Straight Waveguide" sch_x=53 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2207 N$4413 N$4414 "Straight Waveguide" sch_x=53 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2208 N$4415 N$4416 "Straight Waveguide" sch_x=53 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2209 N$4417 N$4418 "Straight Waveguide" sch_x=53 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2210 N$4419 N$4420 "Straight Waveguide" sch_x=53 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2211 N$4421 N$4422 "Straight Waveguide" sch_x=53 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2212 N$4423 N$4424 "Straight Waveguide" sch_x=53 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2213 N$4425 N$4426 "Straight Waveguide" sch_x=53 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2214 N$4427 N$4428 "Straight Waveguide" sch_x=53 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2215 N$4429 N$4430 "Straight Waveguide" sch_x=53 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2216 N$4431 N$4432 "Straight Waveguide" sch_x=53 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2217 N$4433 N$4434 "Straight Waveguide" sch_x=53 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2218 N$4435 N$4436 "Straight Waveguide" sch_x=53 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2219 N$4437 N$4438 "Straight Waveguide" sch_x=53 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2220 N$4439 N$4440 "Straight Waveguide" sch_x=53 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2221 N$4441 N$4442 "Straight Waveguide" sch_x=53 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2222 N$4443 N$4444 "Straight Waveguide" sch_x=53 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2223 N$4445 N$4446 "Straight Waveguide" sch_x=53 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2224 N$4447 N$4448 "Straight Waveguide" sch_x=53 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2225 N$4449 N$4450 "Straight Waveguide" sch_x=53 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2226 N$4451 N$4452 "Straight Waveguide" sch_x=53 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2227 N$4453 N$4454 "Straight Waveguide" sch_x=51 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2228 N$4455 N$4456 "Straight Waveguide" sch_x=51 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2229 N$4457 N$4458 "Straight Waveguide" sch_x=51 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2230 N$4459 N$4460 "Straight Waveguide" sch_x=51 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2231 N$4461 N$4462 "Straight Waveguide" sch_x=51 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2232 N$4463 N$4464 "Straight Waveguide" sch_x=51 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2233 N$4465 N$4466 "Straight Waveguide" sch_x=51 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2234 N$4467 N$4468 "Straight Waveguide" sch_x=51 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2235 N$4469 N$4470 "Straight Waveguide" sch_x=51 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2236 N$4471 N$4472 "Straight Waveguide" sch_x=51 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2237 N$4473 N$4474 "Straight Waveguide" sch_x=51 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2238 N$4475 N$4476 "Straight Waveguide" sch_x=51 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2239 N$4477 N$4478 "Straight Waveguide" sch_x=51 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2240 N$4479 N$4480 "Straight Waveguide" sch_x=51 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2241 N$4481 N$4482 "Straight Waveguide" sch_x=51 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2242 N$4483 N$4484 "Straight Waveguide" sch_x=51 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2243 N$4485 N$4486 "Straight Waveguide" sch_x=51 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2244 N$4487 N$4488 "Straight Waveguide" sch_x=51 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2245 N$4489 N$4490 "Straight Waveguide" sch_x=51 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2246 N$4491 N$4492 "Straight Waveguide" sch_x=51 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2247 N$4493 N$4494 "Straight Waveguide" sch_x=49 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2248 N$4495 N$4496 "Straight Waveguide" sch_x=49 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2249 N$4497 N$4498 "Straight Waveguide" sch_x=49 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2250 N$4499 N$4500 "Straight Waveguide" sch_x=49 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2251 N$4501 N$4502 "Straight Waveguide" sch_x=49 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2252 N$4503 N$4504 "Straight Waveguide" sch_x=49 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2253 N$4505 N$4506 "Straight Waveguide" sch_x=49 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2254 N$4507 N$4508 "Straight Waveguide" sch_x=49 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2255 N$4509 N$4510 "Straight Waveguide" sch_x=49 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2256 N$4511 N$4512 "Straight Waveguide" sch_x=49 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2257 N$4513 N$4514 "Straight Waveguide" sch_x=49 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2258 N$4515 N$4516 "Straight Waveguide" sch_x=49 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2259 N$4517 N$4518 "Straight Waveguide" sch_x=49 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2260 N$4519 N$4520 "Straight Waveguide" sch_x=49 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2261 N$4521 N$4522 "Straight Waveguide" sch_x=49 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2262 N$4523 N$4524 "Straight Waveguide" sch_x=49 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2263 N$4525 N$4526 "Straight Waveguide" sch_x=49 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2264 N$4527 N$4528 "Straight Waveguide" sch_x=49 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2265 N$4529 N$4530 "Straight Waveguide" sch_x=47 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2266 N$4531 N$4532 "Straight Waveguide" sch_x=47 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2267 N$4533 N$4534 "Straight Waveguide" sch_x=47 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2268 N$4535 N$4536 "Straight Waveguide" sch_x=47 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2269 N$4537 N$4538 "Straight Waveguide" sch_x=47 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2270 N$4539 N$4540 "Straight Waveguide" sch_x=47 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2271 N$4541 N$4542 "Straight Waveguide" sch_x=47 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2272 N$4543 N$4544 "Straight Waveguide" sch_x=47 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2273 N$4545 N$4546 "Straight Waveguide" sch_x=47 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2274 N$4547 N$4548 "Straight Waveguide" sch_x=47 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2275 N$4549 N$4550 "Straight Waveguide" sch_x=47 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2276 N$4551 N$4552 "Straight Waveguide" sch_x=47 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2277 N$4553 N$4554 "Straight Waveguide" sch_x=47 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2278 N$4555 N$4556 "Straight Waveguide" sch_x=47 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2279 N$4557 N$4558 "Straight Waveguide" sch_x=47 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2280 N$4559 N$4560 "Straight Waveguide" sch_x=47 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2281 N$4561 N$4562 "Straight Waveguide" sch_x=45 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2282 N$4563 N$4564 "Straight Waveguide" sch_x=45 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2283 N$4565 N$4566 "Straight Waveguide" sch_x=45 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2284 N$4567 N$4568 "Straight Waveguide" sch_x=45 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2285 N$4569 N$4570 "Straight Waveguide" sch_x=45 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2286 N$4571 N$4572 "Straight Waveguide" sch_x=45 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2287 N$4573 N$4574 "Straight Waveguide" sch_x=45 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2288 N$4575 N$4576 "Straight Waveguide" sch_x=45 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2289 N$4577 N$4578 "Straight Waveguide" sch_x=45 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2290 N$4579 N$4580 "Straight Waveguide" sch_x=45 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2291 N$4581 N$4582 "Straight Waveguide" sch_x=45 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2292 N$4583 N$4584 "Straight Waveguide" sch_x=45 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2293 N$4585 N$4586 "Straight Waveguide" sch_x=45 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2294 N$4587 N$4588 "Straight Waveguide" sch_x=45 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2295 N$4589 N$4590 "Straight Waveguide" sch_x=43 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2296 N$4591 N$4592 "Straight Waveguide" sch_x=43 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2297 N$4593 N$4594 "Straight Waveguide" sch_x=43 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2298 N$4595 N$4596 "Straight Waveguide" sch_x=43 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2299 N$4597 N$4598 "Straight Waveguide" sch_x=43 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2300 N$4599 N$4600 "Straight Waveguide" sch_x=43 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2301 N$4601 N$4602 "Straight Waveguide" sch_x=43 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2302 N$4603 N$4604 "Straight Waveguide" sch_x=43 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2303 N$4605 N$4606 "Straight Waveguide" sch_x=43 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2304 N$4607 N$4608 "Straight Waveguide" sch_x=43 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2305 N$4609 N$4610 "Straight Waveguide" sch_x=43 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2306 N$4611 N$4612 "Straight Waveguide" sch_x=43 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2307 N$4613 N$4614 "Straight Waveguide" sch_x=41 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2308 N$4615 N$4616 "Straight Waveguide" sch_x=41 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2309 N$4617 N$4618 "Straight Waveguide" sch_x=41 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2310 N$4619 N$4620 "Straight Waveguide" sch_x=41 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2311 N$4621 N$4622 "Straight Waveguide" sch_x=41 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2312 N$4623 N$4624 "Straight Waveguide" sch_x=41 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2313 N$4625 N$4626 "Straight Waveguide" sch_x=41 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2314 N$4627 N$4628 "Straight Waveguide" sch_x=41 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2315 N$4629 N$4630 "Straight Waveguide" sch_x=41 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2316 N$4631 N$4632 "Straight Waveguide" sch_x=41 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2317 N$4633 N$4634 "Straight Waveguide" sch_x=39 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2318 N$4635 N$4636 "Straight Waveguide" sch_x=39 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2319 N$4637 N$4638 "Straight Waveguide" sch_x=39 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2320 N$4639 N$4640 "Straight Waveguide" sch_x=39 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2321 N$4641 N$4642 "Straight Waveguide" sch_x=39 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2322 N$4643 N$4644 "Straight Waveguide" sch_x=39 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2323 N$4645 N$4646 "Straight Waveguide" sch_x=39 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2324 N$4647 N$4648 "Straight Waveguide" sch_x=39 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2325 N$4649 N$4650 "Straight Waveguide" sch_x=37 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2326 N$4651 N$4652 "Straight Waveguide" sch_x=37 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2327 N$4653 N$4654 "Straight Waveguide" sch_x=37 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2328 N$4655 N$4656 "Straight Waveguide" sch_x=37 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2329 N$4657 N$4658 "Straight Waveguide" sch_x=37 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2330 N$4659 N$4660 "Straight Waveguide" sch_x=37 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2331 N$4661 N$4662 "Straight Waveguide" sch_x=35 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2332 N$4663 N$4664 "Straight Waveguide" sch_x=35 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2333 N$4665 N$4666 "Straight Waveguide" sch_x=35 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2334 N$4667 N$4668 "Straight Waveguide" sch_x=35 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2335 N$4669 N$4670 "Straight Waveguide" sch_x=33 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2336 N$4671 N$4672 "Straight Waveguide" sch_x=33 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2337 N$4674 N$4673 "Straight Waveguide" sch_x=45 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2338 N$4676 N$4675 "Straight Waveguide" sch_x=44 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2339 N$4678 N$4677 "Straight Waveguide" sch_x=43 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2340 N$4680 N$4679 "Straight Waveguide" sch_x=42 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2341 N$4682 N$4681 "Straight Waveguide" sch_x=41 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2342 N$4684 N$4683 "Straight Waveguide" sch_x=40 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2343 N$4686 N$4685 "Straight Waveguide" sch_x=39 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2344 N$4688 N$4687 "Straight Waveguide" sch_x=38 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2345 N$4690 N$4689 "Straight Waveguide" sch_x=37 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2346 N$4692 N$4691 "Straight Waveguide" sch_x=36 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2347 N$4694 N$4693 "Straight Waveguide" sch_x=35 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2348 N$4696 N$4695 "Straight Waveguide" sch_x=34 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2349 N$4698 N$4697 "Straight Waveguide" sch_x=33 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2350 N$4700 N$4699 "Straight Waveguide" sch_x=32 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2351 N$4702 N$4701 "Straight Waveguide" sch_x=31 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2352 N$4704 N$4703 "Straight Waveguide" sch_x=31 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2353 N$4706 N$4705 "Straight Waveguide" sch_x=32 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2354 N$4708 N$4707 "Straight Waveguide" sch_x=33 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2355 N$4710 N$4709 "Straight Waveguide" sch_x=34 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2356 N$4712 N$4711 "Straight Waveguide" sch_x=35 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2357 N$4714 N$4713 "Straight Waveguide" sch_x=36 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2358 N$4716 N$4715 "Straight Waveguide" sch_x=37 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2359 N$4718 N$4717 "Straight Waveguide" sch_x=38 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2360 N$4720 N$4719 "Straight Waveguide" sch_x=39 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2361 N$4722 N$4721 "Straight Waveguide" sch_x=40 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2362 N$4724 N$4723 "Straight Waveguide" sch_x=41 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2363 N$4726 N$4725 "Straight Waveguide" sch_x=42 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2364 N$4728 N$4727 "Straight Waveguide" sch_x=43 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2365 N$4730 N$4729 "Straight Waveguide" sch_x=44 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2366 N$4732 N$4731 "Straight Waveguide" sch_x=45 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2367 N$4734 N$4733 "Straight Waveguide" sch_x=46 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2368 N$4736 N$4735 "Straight Waveguide" sch_x=46 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2369 N$4738 N$4737 "Straight Waveguide" sch_x=-125 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2370 N$4740 N$4739 "Straight Waveguide" sch_x=-125 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2371 N$4742 N$4741 "Straight Waveguide" sch_x=-125 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2372 N$4744 N$4743 "Straight Waveguide" sch_x=-125 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2373 N$4746 N$4745 "Straight Waveguide" sch_x=-125 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2374 N$4748 N$4747 "Straight Waveguide" sch_x=-125 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2375 N$4750 N$4749 "Straight Waveguide" sch_x=-125 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2376 N$4752 N$4751 "Straight Waveguide" sch_x=-125 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2377 N$4754 N$4753 "Straight Waveguide" sch_x=-125 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2378 N$4756 N$4755 "Straight Waveguide" sch_x=-125 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2379 N$4758 N$4757 "Straight Waveguide" sch_x=-125 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2380 N$4760 N$4759 "Straight Waveguide" sch_x=-125 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2381 N$4762 N$4761 "Straight Waveguide" sch_x=-125 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2382 N$4764 N$4763 "Straight Waveguide" sch_x=-125 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2383 N$4766 N$4765 "Straight Waveguide" sch_x=-125 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2384 N$4768 N$4767 "Straight Waveguide" sch_x=-125 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2385 N$4770 N$4769 "Straight Waveguide" sch_x=-125 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2386 N$4772 N$4771 "Straight Waveguide" sch_x=-125 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2387 N$4774 N$4773 "Straight Waveguide" sch_x=-125 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2388 N$4776 N$4775 "Straight Waveguide" sch_x=-125 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2389 N$4778 N$4777 "Straight Waveguide" sch_x=-125 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2390 N$4780 N$4779 "Straight Waveguide" sch_x=-125 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2391 N$4782 N$4781 "Straight Waveguide" sch_x=-125 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2392 N$4784 N$4783 "Straight Waveguide" sch_x=-125 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2393 N$4786 N$4785 "Straight Waveguide" sch_x=-125 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2394 N$4788 N$4787 "Straight Waveguide" sch_x=-125 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2395 N$4790 N$4789 "Straight Waveguide" sch_x=-125 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2396 N$4792 N$4791 "Straight Waveguide" sch_x=-125 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2397 N$4794 N$4793 "Straight Waveguide" sch_x=-125 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2398 N$4796 N$4795 "Straight Waveguide" sch_x=-125 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2399 N$4798 N$4797 "Straight Waveguide" sch_x=-125 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2400 N$4800 N$4799 "Straight Waveguide" sch_x=-125 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2401 N$4802 N$4801 "Straight Waveguide" sch_x=-125 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2402 N$4804 N$4803 "Straight Waveguide" sch_x=-125 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2403 N$4806 N$4805 "Straight Waveguide" sch_x=-125 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2404 N$4808 N$4807 "Straight Waveguide" sch_x=-125 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2405 N$4810 N$4809 "Straight Waveguide" sch_x=-125 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2406 N$4812 N$4811 "Straight Waveguide" sch_x=-125 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2407 N$4814 N$4813 "Straight Waveguide" sch_x=-125 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2408 N$4816 N$4815 "Straight Waveguide" sch_x=-125 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2409 N$4818 N$4817 "Straight Waveguide" sch_x=-125 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2410 N$4820 N$4819 "Straight Waveguide" sch_x=-125 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2411 N$4822 N$4821 "Straight Waveguide" sch_x=-125 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2412 N$4824 N$4823 "Straight Waveguide" sch_x=-125 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2413 N$4826 N$4825 "Straight Waveguide" sch_x=-125 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2414 N$4828 N$4827 "Straight Waveguide" sch_x=-125 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2415 N$4830 N$4829 "Straight Waveguide" sch_x=-125 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2416 N$4832 N$4831 "Straight Waveguide" sch_x=-125 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2417 N$4834 N$4833 "Straight Waveguide" sch_x=-125 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2418 N$4836 N$4835 "Straight Waveguide" sch_x=-125 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2419 N$4838 N$4837 "Straight Waveguide" sch_x=-125 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2420 N$4840 N$4839 "Straight Waveguide" sch_x=-125 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2421 N$4842 N$4841 "Straight Waveguide" sch_x=-125 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2422 N$4844 N$4843 "Straight Waveguide" sch_x=-125 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2423 N$4846 N$4845 "Straight Waveguide" sch_x=-125 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2424 N$4848 N$4847 "Straight Waveguide" sch_x=-125 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2425 N$4850 N$4849 "Straight Waveguide" sch_x=-125 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2426 N$4852 N$4851 "Straight Waveguide" sch_x=-125 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2427 N$4854 N$4853 "Straight Waveguide" sch_x=-125 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2428 N$4856 N$4855 "Straight Waveguide" sch_x=-125 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2429 N$4858 N$4857 "Straight Waveguide" sch_x=-125 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2430 N$4860 N$4859 "Straight Waveguide" sch_x=-125 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2431 N$4862 N$4861 "Straight Waveguide" sch_x=-123 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2432 N$4864 N$4863 "Straight Waveguide" sch_x=-123 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2433 N$4866 N$4865 "Straight Waveguide" sch_x=-123 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2434 N$4868 N$4867 "Straight Waveguide" sch_x=-123 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2435 N$4870 N$4869 "Straight Waveguide" sch_x=-123 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2436 N$4872 N$4871 "Straight Waveguide" sch_x=-123 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2437 N$4874 N$4873 "Straight Waveguide" sch_x=-123 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2438 N$4876 N$4875 "Straight Waveguide" sch_x=-123 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2439 N$4878 N$4877 "Straight Waveguide" sch_x=-123 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2440 N$4880 N$4879 "Straight Waveguide" sch_x=-123 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2441 N$4882 N$4881 "Straight Waveguide" sch_x=-123 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2442 N$4884 N$4883 "Straight Waveguide" sch_x=-123 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2443 N$4886 N$4885 "Straight Waveguide" sch_x=-123 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2444 N$4888 N$4887 "Straight Waveguide" sch_x=-123 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2445 N$4890 N$4889 "Straight Waveguide" sch_x=-123 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2446 N$4892 N$4891 "Straight Waveguide" sch_x=-123 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2447 N$4894 N$4893 "Straight Waveguide" sch_x=-123 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2448 N$4896 N$4895 "Straight Waveguide" sch_x=-123 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2449 N$4898 N$4897 "Straight Waveguide" sch_x=-123 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2450 N$4900 N$4899 "Straight Waveguide" sch_x=-123 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2451 N$4902 N$4901 "Straight Waveguide" sch_x=-123 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2452 N$4904 N$4903 "Straight Waveguide" sch_x=-123 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2453 N$4906 N$4905 "Straight Waveguide" sch_x=-123 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2454 N$4908 N$4907 "Straight Waveguide" sch_x=-123 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2455 N$4910 N$4909 "Straight Waveguide" sch_x=-123 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2456 N$4912 N$4911 "Straight Waveguide" sch_x=-123 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2457 N$4914 N$4913 "Straight Waveguide" sch_x=-123 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2458 N$4916 N$4915 "Straight Waveguide" sch_x=-123 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2459 N$4918 N$4917 "Straight Waveguide" sch_x=-123 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2460 N$4920 N$4919 "Straight Waveguide" sch_x=-123 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2461 N$4922 N$4921 "Straight Waveguide" sch_x=-123 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2462 N$4924 N$4923 "Straight Waveguide" sch_x=-123 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2463 N$4926 N$4925 "Straight Waveguide" sch_x=-123 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2464 N$4928 N$4927 "Straight Waveguide" sch_x=-123 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2465 N$4930 N$4929 "Straight Waveguide" sch_x=-123 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2466 N$4932 N$4931 "Straight Waveguide" sch_x=-123 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2467 N$4934 N$4933 "Straight Waveguide" sch_x=-123 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2468 N$4936 N$4935 "Straight Waveguide" sch_x=-123 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2469 N$4938 N$4937 "Straight Waveguide" sch_x=-123 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2470 N$4940 N$4939 "Straight Waveguide" sch_x=-123 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2471 N$4942 N$4941 "Straight Waveguide" sch_x=-123 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2472 N$4944 N$4943 "Straight Waveguide" sch_x=-123 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2473 N$4946 N$4945 "Straight Waveguide" sch_x=-123 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2474 N$4948 N$4947 "Straight Waveguide" sch_x=-123 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2475 N$4950 N$4949 "Straight Waveguide" sch_x=-123 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2476 N$4952 N$4951 "Straight Waveguide" sch_x=-123 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2477 N$4954 N$4953 "Straight Waveguide" sch_x=-123 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2478 N$4956 N$4955 "Straight Waveguide" sch_x=-123 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2479 N$4958 N$4957 "Straight Waveguide" sch_x=-123 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2480 N$4960 N$4959 "Straight Waveguide" sch_x=-123 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2481 N$4962 N$4961 "Straight Waveguide" sch_x=-123 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2482 N$4964 N$4963 "Straight Waveguide" sch_x=-123 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2483 N$4966 N$4965 "Straight Waveguide" sch_x=-123 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2484 N$4968 N$4967 "Straight Waveguide" sch_x=-123 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2485 N$4970 N$4969 "Straight Waveguide" sch_x=-123 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2486 N$4972 N$4971 "Straight Waveguide" sch_x=-123 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2487 N$4974 N$4973 "Straight Waveguide" sch_x=-123 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2488 N$4976 N$4975 "Straight Waveguide" sch_x=-123 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2489 N$4978 N$4977 "Straight Waveguide" sch_x=-123 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2490 N$4980 N$4979 "Straight Waveguide" sch_x=-123 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2491 N$4982 N$4981 "Straight Waveguide" sch_x=-121 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2492 N$4984 N$4983 "Straight Waveguide" sch_x=-121 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2493 N$4986 N$4985 "Straight Waveguide" sch_x=-121 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2494 N$4988 N$4987 "Straight Waveguide" sch_x=-121 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2495 N$4990 N$4989 "Straight Waveguide" sch_x=-121 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2496 N$4992 N$4991 "Straight Waveguide" sch_x=-121 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2497 N$4994 N$4993 "Straight Waveguide" sch_x=-121 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2498 N$4996 N$4995 "Straight Waveguide" sch_x=-121 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2499 N$4998 N$4997 "Straight Waveguide" sch_x=-121 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2500 N$5000 N$4999 "Straight Waveguide" sch_x=-121 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2501 N$5002 N$5001 "Straight Waveguide" sch_x=-121 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2502 N$5004 N$5003 "Straight Waveguide" sch_x=-121 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2503 N$5006 N$5005 "Straight Waveguide" sch_x=-121 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2504 N$5008 N$5007 "Straight Waveguide" sch_x=-121 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2505 N$5010 N$5009 "Straight Waveguide" sch_x=-121 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2506 N$5012 N$5011 "Straight Waveguide" sch_x=-121 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2507 N$5014 N$5013 "Straight Waveguide" sch_x=-121 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2508 N$5016 N$5015 "Straight Waveguide" sch_x=-121 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2509 N$5018 N$5017 "Straight Waveguide" sch_x=-121 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2510 N$5020 N$5019 "Straight Waveguide" sch_x=-121 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2511 N$5022 N$5021 "Straight Waveguide" sch_x=-121 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2512 N$5024 N$5023 "Straight Waveguide" sch_x=-121 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2513 N$5026 N$5025 "Straight Waveguide" sch_x=-121 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2514 N$5028 N$5027 "Straight Waveguide" sch_x=-121 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2515 N$5030 N$5029 "Straight Waveguide" sch_x=-121 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2516 N$5032 N$5031 "Straight Waveguide" sch_x=-121 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2517 N$5034 N$5033 "Straight Waveguide" sch_x=-121 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2518 N$5036 N$5035 "Straight Waveguide" sch_x=-121 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2519 N$5038 N$5037 "Straight Waveguide" sch_x=-121 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2520 N$5040 N$5039 "Straight Waveguide" sch_x=-121 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2521 N$5042 N$5041 "Straight Waveguide" sch_x=-121 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2522 N$5044 N$5043 "Straight Waveguide" sch_x=-121 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2523 N$5046 N$5045 "Straight Waveguide" sch_x=-121 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2524 N$5048 N$5047 "Straight Waveguide" sch_x=-121 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2525 N$5050 N$5049 "Straight Waveguide" sch_x=-121 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2526 N$5052 N$5051 "Straight Waveguide" sch_x=-121 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2527 N$5054 N$5053 "Straight Waveguide" sch_x=-121 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2528 N$5056 N$5055 "Straight Waveguide" sch_x=-121 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2529 N$5058 N$5057 "Straight Waveguide" sch_x=-121 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2530 N$5060 N$5059 "Straight Waveguide" sch_x=-121 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2531 N$5062 N$5061 "Straight Waveguide" sch_x=-121 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2532 N$5064 N$5063 "Straight Waveguide" sch_x=-121 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2533 N$5066 N$5065 "Straight Waveguide" sch_x=-121 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2534 N$5068 N$5067 "Straight Waveguide" sch_x=-121 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2535 N$5070 N$5069 "Straight Waveguide" sch_x=-121 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2536 N$5072 N$5071 "Straight Waveguide" sch_x=-121 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2537 N$5074 N$5073 "Straight Waveguide" sch_x=-121 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2538 N$5076 N$5075 "Straight Waveguide" sch_x=-121 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2539 N$5078 N$5077 "Straight Waveguide" sch_x=-121 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2540 N$5080 N$5079 "Straight Waveguide" sch_x=-121 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2541 N$5082 N$5081 "Straight Waveguide" sch_x=-121 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2542 N$5084 N$5083 "Straight Waveguide" sch_x=-121 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2543 N$5086 N$5085 "Straight Waveguide" sch_x=-121 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2544 N$5088 N$5087 "Straight Waveguide" sch_x=-121 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2545 N$5090 N$5089 "Straight Waveguide" sch_x=-121 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2546 N$5092 N$5091 "Straight Waveguide" sch_x=-121 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2547 N$5094 N$5093 "Straight Waveguide" sch_x=-121 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2548 N$5096 N$5095 "Straight Waveguide" sch_x=-121 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2549 N$5098 N$5097 "Straight Waveguide" sch_x=-119 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2550 N$5100 N$5099 "Straight Waveguide" sch_x=-119 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2551 N$5102 N$5101 "Straight Waveguide" sch_x=-119 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2552 N$5104 N$5103 "Straight Waveguide" sch_x=-119 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2553 N$5106 N$5105 "Straight Waveguide" sch_x=-119 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2554 N$5108 N$5107 "Straight Waveguide" sch_x=-119 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2555 N$5110 N$5109 "Straight Waveguide" sch_x=-119 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2556 N$5112 N$5111 "Straight Waveguide" sch_x=-119 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2557 N$5114 N$5113 "Straight Waveguide" sch_x=-119 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2558 N$5116 N$5115 "Straight Waveguide" sch_x=-119 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2559 N$5118 N$5117 "Straight Waveguide" sch_x=-119 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2560 N$5120 N$5119 "Straight Waveguide" sch_x=-119 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2561 N$5122 N$5121 "Straight Waveguide" sch_x=-119 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2562 N$5124 N$5123 "Straight Waveguide" sch_x=-119 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2563 N$5126 N$5125 "Straight Waveguide" sch_x=-119 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2564 N$5128 N$5127 "Straight Waveguide" sch_x=-119 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2565 N$5130 N$5129 "Straight Waveguide" sch_x=-119 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2566 N$5132 N$5131 "Straight Waveguide" sch_x=-119 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2567 N$5134 N$5133 "Straight Waveguide" sch_x=-119 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2568 N$5136 N$5135 "Straight Waveguide" sch_x=-119 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2569 N$5138 N$5137 "Straight Waveguide" sch_x=-119 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2570 N$5140 N$5139 "Straight Waveguide" sch_x=-119 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2571 N$5142 N$5141 "Straight Waveguide" sch_x=-119 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2572 N$5144 N$5143 "Straight Waveguide" sch_x=-119 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2573 N$5146 N$5145 "Straight Waveguide" sch_x=-119 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2574 N$5148 N$5147 "Straight Waveguide" sch_x=-119 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2575 N$5150 N$5149 "Straight Waveguide" sch_x=-119 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2576 N$5152 N$5151 "Straight Waveguide" sch_x=-119 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2577 N$5154 N$5153 "Straight Waveguide" sch_x=-119 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2578 N$5156 N$5155 "Straight Waveguide" sch_x=-119 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2579 N$5158 N$5157 "Straight Waveguide" sch_x=-119 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2580 N$5160 N$5159 "Straight Waveguide" sch_x=-119 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2581 N$5162 N$5161 "Straight Waveguide" sch_x=-119 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2582 N$5164 N$5163 "Straight Waveguide" sch_x=-119 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2583 N$5166 N$5165 "Straight Waveguide" sch_x=-119 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2584 N$5168 N$5167 "Straight Waveguide" sch_x=-119 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2585 N$5170 N$5169 "Straight Waveguide" sch_x=-119 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2586 N$5172 N$5171 "Straight Waveguide" sch_x=-119 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2587 N$5174 N$5173 "Straight Waveguide" sch_x=-119 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2588 N$5176 N$5175 "Straight Waveguide" sch_x=-119 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2589 N$5178 N$5177 "Straight Waveguide" sch_x=-119 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2590 N$5180 N$5179 "Straight Waveguide" sch_x=-119 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2591 N$5182 N$5181 "Straight Waveguide" sch_x=-119 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2592 N$5184 N$5183 "Straight Waveguide" sch_x=-119 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2593 N$5186 N$5185 "Straight Waveguide" sch_x=-119 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2594 N$5188 N$5187 "Straight Waveguide" sch_x=-119 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2595 N$5190 N$5189 "Straight Waveguide" sch_x=-119 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2596 N$5192 N$5191 "Straight Waveguide" sch_x=-119 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2597 N$5194 N$5193 "Straight Waveguide" sch_x=-119 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2598 N$5196 N$5195 "Straight Waveguide" sch_x=-119 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2599 N$5198 N$5197 "Straight Waveguide" sch_x=-119 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2600 N$5200 N$5199 "Straight Waveguide" sch_x=-119 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2601 N$5202 N$5201 "Straight Waveguide" sch_x=-119 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2602 N$5204 N$5203 "Straight Waveguide" sch_x=-119 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2603 N$5206 N$5205 "Straight Waveguide" sch_x=-119 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2604 N$5208 N$5207 "Straight Waveguide" sch_x=-119 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2605 N$5210 N$5209 "Straight Waveguide" sch_x=-117 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2606 N$5212 N$5211 "Straight Waveguide" sch_x=-117 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2607 N$5214 N$5213 "Straight Waveguide" sch_x=-117 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2608 N$5216 N$5215 "Straight Waveguide" sch_x=-117 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2609 N$5218 N$5217 "Straight Waveguide" sch_x=-117 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2610 N$5220 N$5219 "Straight Waveguide" sch_x=-117 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2611 N$5222 N$5221 "Straight Waveguide" sch_x=-117 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2612 N$5224 N$5223 "Straight Waveguide" sch_x=-117 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2613 N$5226 N$5225 "Straight Waveguide" sch_x=-117 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2614 N$5228 N$5227 "Straight Waveguide" sch_x=-117 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2615 N$5230 N$5229 "Straight Waveguide" sch_x=-117 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2616 N$5232 N$5231 "Straight Waveguide" sch_x=-117 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2617 N$5234 N$5233 "Straight Waveguide" sch_x=-117 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2618 N$5236 N$5235 "Straight Waveguide" sch_x=-117 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2619 N$5238 N$5237 "Straight Waveguide" sch_x=-117 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2620 N$5240 N$5239 "Straight Waveguide" sch_x=-117 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2621 N$5242 N$5241 "Straight Waveguide" sch_x=-117 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2622 N$5244 N$5243 "Straight Waveguide" sch_x=-117 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2623 N$5246 N$5245 "Straight Waveguide" sch_x=-117 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2624 N$5248 N$5247 "Straight Waveguide" sch_x=-117 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2625 N$5250 N$5249 "Straight Waveguide" sch_x=-117 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2626 N$5252 N$5251 "Straight Waveguide" sch_x=-117 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2627 N$5254 N$5253 "Straight Waveguide" sch_x=-117 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2628 N$5256 N$5255 "Straight Waveguide" sch_x=-117 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2629 N$5258 N$5257 "Straight Waveguide" sch_x=-117 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2630 N$5260 N$5259 "Straight Waveguide" sch_x=-117 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2631 N$5262 N$5261 "Straight Waveguide" sch_x=-117 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2632 N$5264 N$5263 "Straight Waveguide" sch_x=-117 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2633 N$5266 N$5265 "Straight Waveguide" sch_x=-117 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2634 N$5268 N$5267 "Straight Waveguide" sch_x=-117 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2635 N$5270 N$5269 "Straight Waveguide" sch_x=-117 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2636 N$5272 N$5271 "Straight Waveguide" sch_x=-117 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2637 N$5274 N$5273 "Straight Waveguide" sch_x=-117 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2638 N$5276 N$5275 "Straight Waveguide" sch_x=-117 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2639 N$5278 N$5277 "Straight Waveguide" sch_x=-117 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2640 N$5280 N$5279 "Straight Waveguide" sch_x=-117 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2641 N$5282 N$5281 "Straight Waveguide" sch_x=-117 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2642 N$5284 N$5283 "Straight Waveguide" sch_x=-117 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2643 N$5286 N$5285 "Straight Waveguide" sch_x=-117 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2644 N$5288 N$5287 "Straight Waveguide" sch_x=-117 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2645 N$5290 N$5289 "Straight Waveguide" sch_x=-117 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2646 N$5292 N$5291 "Straight Waveguide" sch_x=-117 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2647 N$5294 N$5293 "Straight Waveguide" sch_x=-117 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2648 N$5296 N$5295 "Straight Waveguide" sch_x=-117 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2649 N$5298 N$5297 "Straight Waveguide" sch_x=-117 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2650 N$5300 N$5299 "Straight Waveguide" sch_x=-117 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2651 N$5302 N$5301 "Straight Waveguide" sch_x=-117 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2652 N$5304 N$5303 "Straight Waveguide" sch_x=-117 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2653 N$5306 N$5305 "Straight Waveguide" sch_x=-117 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2654 N$5308 N$5307 "Straight Waveguide" sch_x=-117 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2655 N$5310 N$5309 "Straight Waveguide" sch_x=-117 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2656 N$5312 N$5311 "Straight Waveguide" sch_x=-117 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2657 N$5314 N$5313 "Straight Waveguide" sch_x=-117 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2658 N$5316 N$5315 "Straight Waveguide" sch_x=-117 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2659 N$5318 N$5317 "Straight Waveguide" sch_x=-115 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2660 N$5320 N$5319 "Straight Waveguide" sch_x=-115 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2661 N$5322 N$5321 "Straight Waveguide" sch_x=-115 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2662 N$5324 N$5323 "Straight Waveguide" sch_x=-115 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2663 N$5326 N$5325 "Straight Waveguide" sch_x=-115 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2664 N$5328 N$5327 "Straight Waveguide" sch_x=-115 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2665 N$5330 N$5329 "Straight Waveguide" sch_x=-115 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2666 N$5332 N$5331 "Straight Waveguide" sch_x=-115 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2667 N$5334 N$5333 "Straight Waveguide" sch_x=-115 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2668 N$5336 N$5335 "Straight Waveguide" sch_x=-115 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2669 N$5338 N$5337 "Straight Waveguide" sch_x=-115 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2670 N$5340 N$5339 "Straight Waveguide" sch_x=-115 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2671 N$5342 N$5341 "Straight Waveguide" sch_x=-115 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2672 N$5344 N$5343 "Straight Waveguide" sch_x=-115 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2673 N$5346 N$5345 "Straight Waveguide" sch_x=-115 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2674 N$5348 N$5347 "Straight Waveguide" sch_x=-115 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2675 N$5350 N$5349 "Straight Waveguide" sch_x=-115 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2676 N$5352 N$5351 "Straight Waveguide" sch_x=-115 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2677 N$5354 N$5353 "Straight Waveguide" sch_x=-115 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2678 N$5356 N$5355 "Straight Waveguide" sch_x=-115 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2679 N$5358 N$5357 "Straight Waveguide" sch_x=-115 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2680 N$5360 N$5359 "Straight Waveguide" sch_x=-115 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2681 N$5362 N$5361 "Straight Waveguide" sch_x=-115 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2682 N$5364 N$5363 "Straight Waveguide" sch_x=-115 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2683 N$5366 N$5365 "Straight Waveguide" sch_x=-115 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2684 N$5368 N$5367 "Straight Waveguide" sch_x=-115 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2685 N$5370 N$5369 "Straight Waveguide" sch_x=-115 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2686 N$5372 N$5371 "Straight Waveguide" sch_x=-115 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2687 N$5374 N$5373 "Straight Waveguide" sch_x=-115 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2688 N$5376 N$5375 "Straight Waveguide" sch_x=-115 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2689 N$5378 N$5377 "Straight Waveguide" sch_x=-115 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2690 N$5380 N$5379 "Straight Waveguide" sch_x=-115 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2691 N$5382 N$5381 "Straight Waveguide" sch_x=-115 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2692 N$5384 N$5383 "Straight Waveguide" sch_x=-115 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2693 N$5386 N$5385 "Straight Waveguide" sch_x=-115 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2694 N$5388 N$5387 "Straight Waveguide" sch_x=-115 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2695 N$5390 N$5389 "Straight Waveguide" sch_x=-115 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2696 N$5392 N$5391 "Straight Waveguide" sch_x=-115 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2697 N$5394 N$5393 "Straight Waveguide" sch_x=-115 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2698 N$5396 N$5395 "Straight Waveguide" sch_x=-115 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2699 N$5398 N$5397 "Straight Waveguide" sch_x=-115 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2700 N$5400 N$5399 "Straight Waveguide" sch_x=-115 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2701 N$5402 N$5401 "Straight Waveguide" sch_x=-115 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2702 N$5404 N$5403 "Straight Waveguide" sch_x=-115 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2703 N$5406 N$5405 "Straight Waveguide" sch_x=-115 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2704 N$5408 N$5407 "Straight Waveguide" sch_x=-115 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2705 N$5410 N$5409 "Straight Waveguide" sch_x=-115 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2706 N$5412 N$5411 "Straight Waveguide" sch_x=-115 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2707 N$5414 N$5413 "Straight Waveguide" sch_x=-115 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2708 N$5416 N$5415 "Straight Waveguide" sch_x=-115 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2709 N$5418 N$5417 "Straight Waveguide" sch_x=-115 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2710 N$5420 N$5419 "Straight Waveguide" sch_x=-115 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2711 N$5422 N$5421 "Straight Waveguide" sch_x=-113 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2712 N$5424 N$5423 "Straight Waveguide" sch_x=-113 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2713 N$5426 N$5425 "Straight Waveguide" sch_x=-113 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2714 N$5428 N$5427 "Straight Waveguide" sch_x=-113 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2715 N$5430 N$5429 "Straight Waveguide" sch_x=-113 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2716 N$5432 N$5431 "Straight Waveguide" sch_x=-113 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2717 N$5434 N$5433 "Straight Waveguide" sch_x=-113 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2718 N$5436 N$5435 "Straight Waveguide" sch_x=-113 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2719 N$5438 N$5437 "Straight Waveguide" sch_x=-113 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2720 N$5440 N$5439 "Straight Waveguide" sch_x=-113 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2721 N$5442 N$5441 "Straight Waveguide" sch_x=-113 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2722 N$5444 N$5443 "Straight Waveguide" sch_x=-113 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2723 N$5446 N$5445 "Straight Waveguide" sch_x=-113 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2724 N$5448 N$5447 "Straight Waveguide" sch_x=-113 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2725 N$5450 N$5449 "Straight Waveguide" sch_x=-113 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2726 N$5452 N$5451 "Straight Waveguide" sch_x=-113 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2727 N$5454 N$5453 "Straight Waveguide" sch_x=-113 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2728 N$5456 N$5455 "Straight Waveguide" sch_x=-113 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2729 N$5458 N$5457 "Straight Waveguide" sch_x=-113 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2730 N$5460 N$5459 "Straight Waveguide" sch_x=-113 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2731 N$5462 N$5461 "Straight Waveguide" sch_x=-113 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2732 N$5464 N$5463 "Straight Waveguide" sch_x=-113 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2733 N$5466 N$5465 "Straight Waveguide" sch_x=-113 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2734 N$5468 N$5467 "Straight Waveguide" sch_x=-113 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2735 N$5470 N$5469 "Straight Waveguide" sch_x=-113 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2736 N$5472 N$5471 "Straight Waveguide" sch_x=-113 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2737 N$5474 N$5473 "Straight Waveguide" sch_x=-113 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2738 N$5476 N$5475 "Straight Waveguide" sch_x=-113 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2739 N$5478 N$5477 "Straight Waveguide" sch_x=-113 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2740 N$5480 N$5479 "Straight Waveguide" sch_x=-113 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2741 N$5482 N$5481 "Straight Waveguide" sch_x=-113 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2742 N$5484 N$5483 "Straight Waveguide" sch_x=-113 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2743 N$5486 N$5485 "Straight Waveguide" sch_x=-113 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2744 N$5488 N$5487 "Straight Waveguide" sch_x=-113 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2745 N$5490 N$5489 "Straight Waveguide" sch_x=-113 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2746 N$5492 N$5491 "Straight Waveguide" sch_x=-113 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2747 N$5494 N$5493 "Straight Waveguide" sch_x=-113 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2748 N$5496 N$5495 "Straight Waveguide" sch_x=-113 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2749 N$5498 N$5497 "Straight Waveguide" sch_x=-113 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2750 N$5500 N$5499 "Straight Waveguide" sch_x=-113 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2751 N$5502 N$5501 "Straight Waveguide" sch_x=-113 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2752 N$5504 N$5503 "Straight Waveguide" sch_x=-113 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2753 N$5506 N$5505 "Straight Waveguide" sch_x=-113 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2754 N$5508 N$5507 "Straight Waveguide" sch_x=-113 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2755 N$5510 N$5509 "Straight Waveguide" sch_x=-113 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2756 N$5512 N$5511 "Straight Waveguide" sch_x=-113 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2757 N$5514 N$5513 "Straight Waveguide" sch_x=-113 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2758 N$5516 N$5515 "Straight Waveguide" sch_x=-113 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2759 N$5518 N$5517 "Straight Waveguide" sch_x=-113 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2760 N$5520 N$5519 "Straight Waveguide" sch_x=-113 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2761 N$5522 N$5521 "Straight Waveguide" sch_x=-111 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2762 N$5524 N$5523 "Straight Waveguide" sch_x=-111 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2763 N$5526 N$5525 "Straight Waveguide" sch_x=-111 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2764 N$5528 N$5527 "Straight Waveguide" sch_x=-111 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2765 N$5530 N$5529 "Straight Waveguide" sch_x=-111 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2766 N$5532 N$5531 "Straight Waveguide" sch_x=-111 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2767 N$5534 N$5533 "Straight Waveguide" sch_x=-111 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2768 N$5536 N$5535 "Straight Waveguide" sch_x=-111 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2769 N$5538 N$5537 "Straight Waveguide" sch_x=-111 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2770 N$5540 N$5539 "Straight Waveguide" sch_x=-111 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2771 N$5542 N$5541 "Straight Waveguide" sch_x=-111 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2772 N$5544 N$5543 "Straight Waveguide" sch_x=-111 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2773 N$5546 N$5545 "Straight Waveguide" sch_x=-111 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2774 N$5548 N$5547 "Straight Waveguide" sch_x=-111 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2775 N$5550 N$5549 "Straight Waveguide" sch_x=-111 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2776 N$5552 N$5551 "Straight Waveguide" sch_x=-111 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2777 N$5554 N$5553 "Straight Waveguide" sch_x=-111 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2778 N$5556 N$5555 "Straight Waveguide" sch_x=-111 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2779 N$5558 N$5557 "Straight Waveguide" sch_x=-111 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2780 N$5560 N$5559 "Straight Waveguide" sch_x=-111 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2781 N$5562 N$5561 "Straight Waveguide" sch_x=-111 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2782 N$5564 N$5563 "Straight Waveguide" sch_x=-111 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2783 N$5566 N$5565 "Straight Waveguide" sch_x=-111 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2784 N$5568 N$5567 "Straight Waveguide" sch_x=-111 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2785 N$5570 N$5569 "Straight Waveguide" sch_x=-111 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2786 N$5572 N$5571 "Straight Waveguide" sch_x=-111 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2787 N$5574 N$5573 "Straight Waveguide" sch_x=-111 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2788 N$5576 N$5575 "Straight Waveguide" sch_x=-111 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2789 N$5578 N$5577 "Straight Waveguide" sch_x=-111 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2790 N$5580 N$5579 "Straight Waveguide" sch_x=-111 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2791 N$5582 N$5581 "Straight Waveguide" sch_x=-111 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2792 N$5584 N$5583 "Straight Waveguide" sch_x=-111 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2793 N$5586 N$5585 "Straight Waveguide" sch_x=-111 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2794 N$5588 N$5587 "Straight Waveguide" sch_x=-111 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2795 N$5590 N$5589 "Straight Waveguide" sch_x=-111 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2796 N$5592 N$5591 "Straight Waveguide" sch_x=-111 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2797 N$5594 N$5593 "Straight Waveguide" sch_x=-111 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2798 N$5596 N$5595 "Straight Waveguide" sch_x=-111 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2799 N$5598 N$5597 "Straight Waveguide" sch_x=-111 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2800 N$5600 N$5599 "Straight Waveguide" sch_x=-111 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2801 N$5602 N$5601 "Straight Waveguide" sch_x=-111 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2802 N$5604 N$5603 "Straight Waveguide" sch_x=-111 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2803 N$5606 N$5605 "Straight Waveguide" sch_x=-111 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2804 N$5608 N$5607 "Straight Waveguide" sch_x=-111 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2805 N$5610 N$5609 "Straight Waveguide" sch_x=-111 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2806 N$5612 N$5611 "Straight Waveguide" sch_x=-111 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2807 N$5614 N$5613 "Straight Waveguide" sch_x=-111 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2808 N$5616 N$5615 "Straight Waveguide" sch_x=-111 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2809 N$5618 N$5617 "Straight Waveguide" sch_x=-109 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2810 N$5620 N$5619 "Straight Waveguide" sch_x=-109 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2811 N$5622 N$5621 "Straight Waveguide" sch_x=-109 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2812 N$5624 N$5623 "Straight Waveguide" sch_x=-109 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2813 N$5626 N$5625 "Straight Waveguide" sch_x=-109 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2814 N$5628 N$5627 "Straight Waveguide" sch_x=-109 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2815 N$5630 N$5629 "Straight Waveguide" sch_x=-109 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2816 N$5632 N$5631 "Straight Waveguide" sch_x=-109 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2817 N$5634 N$5633 "Straight Waveguide" sch_x=-109 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2818 N$5636 N$5635 "Straight Waveguide" sch_x=-109 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2819 N$5638 N$5637 "Straight Waveguide" sch_x=-109 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2820 N$5640 N$5639 "Straight Waveguide" sch_x=-109 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2821 N$5642 N$5641 "Straight Waveguide" sch_x=-109 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2822 N$5644 N$5643 "Straight Waveguide" sch_x=-109 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2823 N$5646 N$5645 "Straight Waveguide" sch_x=-109 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2824 N$5648 N$5647 "Straight Waveguide" sch_x=-109 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2825 N$5650 N$5649 "Straight Waveguide" sch_x=-109 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2826 N$5652 N$5651 "Straight Waveguide" sch_x=-109 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2827 N$5654 N$5653 "Straight Waveguide" sch_x=-109 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2828 N$5656 N$5655 "Straight Waveguide" sch_x=-109 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2829 N$5658 N$5657 "Straight Waveguide" sch_x=-109 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2830 N$5660 N$5659 "Straight Waveguide" sch_x=-109 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2831 N$5662 N$5661 "Straight Waveguide" sch_x=-109 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2832 N$5664 N$5663 "Straight Waveguide" sch_x=-109 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2833 N$5666 N$5665 "Straight Waveguide" sch_x=-109 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2834 N$5668 N$5667 "Straight Waveguide" sch_x=-109 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2835 N$5670 N$5669 "Straight Waveguide" sch_x=-109 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2836 N$5672 N$5671 "Straight Waveguide" sch_x=-109 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2837 N$5674 N$5673 "Straight Waveguide" sch_x=-109 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2838 N$5676 N$5675 "Straight Waveguide" sch_x=-109 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2839 N$5678 N$5677 "Straight Waveguide" sch_x=-109 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2840 N$5680 N$5679 "Straight Waveguide" sch_x=-109 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2841 N$5682 N$5681 "Straight Waveguide" sch_x=-109 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2842 N$5684 N$5683 "Straight Waveguide" sch_x=-109 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2843 N$5686 N$5685 "Straight Waveguide" sch_x=-109 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2844 N$5688 N$5687 "Straight Waveguide" sch_x=-109 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2845 N$5690 N$5689 "Straight Waveguide" sch_x=-109 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2846 N$5692 N$5691 "Straight Waveguide" sch_x=-109 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2847 N$5694 N$5693 "Straight Waveguide" sch_x=-109 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2848 N$5696 N$5695 "Straight Waveguide" sch_x=-109 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2849 N$5698 N$5697 "Straight Waveguide" sch_x=-109 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2850 N$5700 N$5699 "Straight Waveguide" sch_x=-109 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2851 N$5702 N$5701 "Straight Waveguide" sch_x=-109 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2852 N$5704 N$5703 "Straight Waveguide" sch_x=-109 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2853 N$5706 N$5705 "Straight Waveguide" sch_x=-109 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2854 N$5708 N$5707 "Straight Waveguide" sch_x=-109 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2855 N$5710 N$5709 "Straight Waveguide" sch_x=-107 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2856 N$5712 N$5711 "Straight Waveguide" sch_x=-107 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2857 N$5714 N$5713 "Straight Waveguide" sch_x=-107 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2858 N$5716 N$5715 "Straight Waveguide" sch_x=-107 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2859 N$5718 N$5717 "Straight Waveguide" sch_x=-107 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2860 N$5720 N$5719 "Straight Waveguide" sch_x=-107 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2861 N$5722 N$5721 "Straight Waveguide" sch_x=-107 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2862 N$5724 N$5723 "Straight Waveguide" sch_x=-107 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2863 N$5726 N$5725 "Straight Waveguide" sch_x=-107 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2864 N$5728 N$5727 "Straight Waveguide" sch_x=-107 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2865 N$5730 N$5729 "Straight Waveguide" sch_x=-107 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2866 N$5732 N$5731 "Straight Waveguide" sch_x=-107 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2867 N$5734 N$5733 "Straight Waveguide" sch_x=-107 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2868 N$5736 N$5735 "Straight Waveguide" sch_x=-107 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2869 N$5738 N$5737 "Straight Waveguide" sch_x=-107 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2870 N$5740 N$5739 "Straight Waveguide" sch_x=-107 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2871 N$5742 N$5741 "Straight Waveguide" sch_x=-107 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2872 N$5744 N$5743 "Straight Waveguide" sch_x=-107 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2873 N$5746 N$5745 "Straight Waveguide" sch_x=-107 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2874 N$5748 N$5747 "Straight Waveguide" sch_x=-107 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2875 N$5750 N$5749 "Straight Waveguide" sch_x=-107 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2876 N$5752 N$5751 "Straight Waveguide" sch_x=-107 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2877 N$5754 N$5753 "Straight Waveguide" sch_x=-107 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2878 N$5756 N$5755 "Straight Waveguide" sch_x=-107 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2879 N$5758 N$5757 "Straight Waveguide" sch_x=-107 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2880 N$5760 N$5759 "Straight Waveguide" sch_x=-107 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2881 N$5762 N$5761 "Straight Waveguide" sch_x=-107 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2882 N$5764 N$5763 "Straight Waveguide" sch_x=-107 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2883 N$5766 N$5765 "Straight Waveguide" sch_x=-107 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2884 N$5768 N$5767 "Straight Waveguide" sch_x=-107 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2885 N$5770 N$5769 "Straight Waveguide" sch_x=-107 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2886 N$5772 N$5771 "Straight Waveguide" sch_x=-107 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2887 N$5774 N$5773 "Straight Waveguide" sch_x=-107 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2888 N$5776 N$5775 "Straight Waveguide" sch_x=-107 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2889 N$5778 N$5777 "Straight Waveguide" sch_x=-107 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2890 N$5780 N$5779 "Straight Waveguide" sch_x=-107 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2891 N$5782 N$5781 "Straight Waveguide" sch_x=-107 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2892 N$5784 N$5783 "Straight Waveguide" sch_x=-107 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2893 N$5786 N$5785 "Straight Waveguide" sch_x=-107 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2894 N$5788 N$5787 "Straight Waveguide" sch_x=-107 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2895 N$5790 N$5789 "Straight Waveguide" sch_x=-107 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2896 N$5792 N$5791 "Straight Waveguide" sch_x=-107 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2897 N$5794 N$5793 "Straight Waveguide" sch_x=-107 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2898 N$5796 N$5795 "Straight Waveguide" sch_x=-107 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2899 N$5798 N$5797 "Straight Waveguide" sch_x=-105 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2900 N$5800 N$5799 "Straight Waveguide" sch_x=-105 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2901 N$5802 N$5801 "Straight Waveguide" sch_x=-105 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2902 N$5804 N$5803 "Straight Waveguide" sch_x=-105 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2903 N$5806 N$5805 "Straight Waveguide" sch_x=-105 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2904 N$5808 N$5807 "Straight Waveguide" sch_x=-105 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2905 N$5810 N$5809 "Straight Waveguide" sch_x=-105 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2906 N$5812 N$5811 "Straight Waveguide" sch_x=-105 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2907 N$5814 N$5813 "Straight Waveguide" sch_x=-105 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2908 N$5816 N$5815 "Straight Waveguide" sch_x=-105 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2909 N$5818 N$5817 "Straight Waveguide" sch_x=-105 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2910 N$5820 N$5819 "Straight Waveguide" sch_x=-105 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2911 N$5822 N$5821 "Straight Waveguide" sch_x=-105 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2912 N$5824 N$5823 "Straight Waveguide" sch_x=-105 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2913 N$5826 N$5825 "Straight Waveguide" sch_x=-105 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2914 N$5828 N$5827 "Straight Waveguide" sch_x=-105 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2915 N$5830 N$5829 "Straight Waveguide" sch_x=-105 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2916 N$5832 N$5831 "Straight Waveguide" sch_x=-105 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2917 N$5834 N$5833 "Straight Waveguide" sch_x=-105 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2918 N$5836 N$5835 "Straight Waveguide" sch_x=-105 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2919 N$5838 N$5837 "Straight Waveguide" sch_x=-105 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2920 N$5840 N$5839 "Straight Waveguide" sch_x=-105 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2921 N$5842 N$5841 "Straight Waveguide" sch_x=-105 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2922 N$5844 N$5843 "Straight Waveguide" sch_x=-105 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2923 N$5846 N$5845 "Straight Waveguide" sch_x=-105 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2924 N$5848 N$5847 "Straight Waveguide" sch_x=-105 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2925 N$5850 N$5849 "Straight Waveguide" sch_x=-105 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2926 N$5852 N$5851 "Straight Waveguide" sch_x=-105 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2927 N$5854 N$5853 "Straight Waveguide" sch_x=-105 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2928 N$5856 N$5855 "Straight Waveguide" sch_x=-105 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2929 N$5858 N$5857 "Straight Waveguide" sch_x=-105 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2930 N$5860 N$5859 "Straight Waveguide" sch_x=-105 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2931 N$5862 N$5861 "Straight Waveguide" sch_x=-105 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2932 N$5864 N$5863 "Straight Waveguide" sch_x=-105 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2933 N$5866 N$5865 "Straight Waveguide" sch_x=-105 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2934 N$5868 N$5867 "Straight Waveguide" sch_x=-105 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2935 N$5870 N$5869 "Straight Waveguide" sch_x=-105 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2936 N$5872 N$5871 "Straight Waveguide" sch_x=-105 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2937 N$5874 N$5873 "Straight Waveguide" sch_x=-105 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2938 N$5876 N$5875 "Straight Waveguide" sch_x=-105 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2939 N$5878 N$5877 "Straight Waveguide" sch_x=-105 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2940 N$5880 N$5879 "Straight Waveguide" sch_x=-105 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2941 N$5882 N$5881 "Straight Waveguide" sch_x=-103 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2942 N$5884 N$5883 "Straight Waveguide" sch_x=-103 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2943 N$5886 N$5885 "Straight Waveguide" sch_x=-103 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2944 N$5888 N$5887 "Straight Waveguide" sch_x=-103 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2945 N$5890 N$5889 "Straight Waveguide" sch_x=-103 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2946 N$5892 N$5891 "Straight Waveguide" sch_x=-103 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2947 N$5894 N$5893 "Straight Waveguide" sch_x=-103 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2948 N$5896 N$5895 "Straight Waveguide" sch_x=-103 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2949 N$5898 N$5897 "Straight Waveguide" sch_x=-103 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2950 N$5900 N$5899 "Straight Waveguide" sch_x=-103 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2951 N$5902 N$5901 "Straight Waveguide" sch_x=-103 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2952 N$5904 N$5903 "Straight Waveguide" sch_x=-103 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2953 N$5906 N$5905 "Straight Waveguide" sch_x=-103 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2954 N$5908 N$5907 "Straight Waveguide" sch_x=-103 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2955 N$5910 N$5909 "Straight Waveguide" sch_x=-103 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2956 N$5912 N$5911 "Straight Waveguide" sch_x=-103 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2957 N$5914 N$5913 "Straight Waveguide" sch_x=-103 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2958 N$5916 N$5915 "Straight Waveguide" sch_x=-103 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2959 N$5918 N$5917 "Straight Waveguide" sch_x=-103 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2960 N$5920 N$5919 "Straight Waveguide" sch_x=-103 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2961 N$5922 N$5921 "Straight Waveguide" sch_x=-103 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2962 N$5924 N$5923 "Straight Waveguide" sch_x=-103 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2963 N$5926 N$5925 "Straight Waveguide" sch_x=-103 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2964 N$5928 N$5927 "Straight Waveguide" sch_x=-103 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2965 N$5930 N$5929 "Straight Waveguide" sch_x=-103 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2966 N$5932 N$5931 "Straight Waveguide" sch_x=-103 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2967 N$5934 N$5933 "Straight Waveguide" sch_x=-103 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2968 N$5936 N$5935 "Straight Waveguide" sch_x=-103 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2969 N$5938 N$5937 "Straight Waveguide" sch_x=-103 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2970 N$5940 N$5939 "Straight Waveguide" sch_x=-103 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2971 N$5942 N$5941 "Straight Waveguide" sch_x=-103 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2972 N$5944 N$5943 "Straight Waveguide" sch_x=-103 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2973 N$5946 N$5945 "Straight Waveguide" sch_x=-103 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2974 N$5948 N$5947 "Straight Waveguide" sch_x=-103 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2975 N$5950 N$5949 "Straight Waveguide" sch_x=-103 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2976 N$5952 N$5951 "Straight Waveguide" sch_x=-103 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2977 N$5954 N$5953 "Straight Waveguide" sch_x=-103 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2978 N$5956 N$5955 "Straight Waveguide" sch_x=-103 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2979 N$5958 N$5957 "Straight Waveguide" sch_x=-103 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2980 N$5960 N$5959 "Straight Waveguide" sch_x=-103 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2981 N$5962 N$5961 "Straight Waveguide" sch_x=-101 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2982 N$5964 N$5963 "Straight Waveguide" sch_x=-101 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2983 N$5966 N$5965 "Straight Waveguide" sch_x=-101 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2984 N$5968 N$5967 "Straight Waveguide" sch_x=-101 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2985 N$5970 N$5969 "Straight Waveguide" sch_x=-101 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2986 N$5972 N$5971 "Straight Waveguide" sch_x=-101 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2987 N$5974 N$5973 "Straight Waveguide" sch_x=-101 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2988 N$5976 N$5975 "Straight Waveguide" sch_x=-101 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2989 N$5978 N$5977 "Straight Waveguide" sch_x=-101 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2990 N$5980 N$5979 "Straight Waveguide" sch_x=-101 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2991 N$5982 N$5981 "Straight Waveguide" sch_x=-101 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2992 N$5984 N$5983 "Straight Waveguide" sch_x=-101 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2993 N$5986 N$5985 "Straight Waveguide" sch_x=-101 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2994 N$5988 N$5987 "Straight Waveguide" sch_x=-101 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2995 N$5990 N$5989 "Straight Waveguide" sch_x=-101 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2996 N$5992 N$5991 "Straight Waveguide" sch_x=-101 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2997 N$5994 N$5993 "Straight Waveguide" sch_x=-101 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2998 N$5996 N$5995 "Straight Waveguide" sch_x=-101 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2999 N$5998 N$5997 "Straight Waveguide" sch_x=-101 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3000 N$6000 N$5999 "Straight Waveguide" sch_x=-101 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3001 N$6002 N$6001 "Straight Waveguide" sch_x=-101 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3002 N$6004 N$6003 "Straight Waveguide" sch_x=-101 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3003 N$6006 N$6005 "Straight Waveguide" sch_x=-101 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3004 N$6008 N$6007 "Straight Waveguide" sch_x=-101 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3005 N$6010 N$6009 "Straight Waveguide" sch_x=-101 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3006 N$6012 N$6011 "Straight Waveguide" sch_x=-101 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3007 N$6014 N$6013 "Straight Waveguide" sch_x=-101 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3008 N$6016 N$6015 "Straight Waveguide" sch_x=-101 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3009 N$6018 N$6017 "Straight Waveguide" sch_x=-101 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3010 N$6020 N$6019 "Straight Waveguide" sch_x=-101 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3011 N$6022 N$6021 "Straight Waveguide" sch_x=-101 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3012 N$6024 N$6023 "Straight Waveguide" sch_x=-101 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3013 N$6026 N$6025 "Straight Waveguide" sch_x=-101 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3014 N$6028 N$6027 "Straight Waveguide" sch_x=-101 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3015 N$6030 N$6029 "Straight Waveguide" sch_x=-101 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3016 N$6032 N$6031 "Straight Waveguide" sch_x=-101 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3017 N$6034 N$6033 "Straight Waveguide" sch_x=-101 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3018 N$6036 N$6035 "Straight Waveguide" sch_x=-101 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3019 N$6038 N$6037 "Straight Waveguide" sch_x=-99 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3020 N$6040 N$6039 "Straight Waveguide" sch_x=-99 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3021 N$6042 N$6041 "Straight Waveguide" sch_x=-99 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3022 N$6044 N$6043 "Straight Waveguide" sch_x=-99 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3023 N$6046 N$6045 "Straight Waveguide" sch_x=-99 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3024 N$6048 N$6047 "Straight Waveguide" sch_x=-99 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3025 N$6050 N$6049 "Straight Waveguide" sch_x=-99 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3026 N$6052 N$6051 "Straight Waveguide" sch_x=-99 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3027 N$6054 N$6053 "Straight Waveguide" sch_x=-99 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3028 N$6056 N$6055 "Straight Waveguide" sch_x=-99 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3029 N$6058 N$6057 "Straight Waveguide" sch_x=-99 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3030 N$6060 N$6059 "Straight Waveguide" sch_x=-99 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3031 N$6062 N$6061 "Straight Waveguide" sch_x=-99 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3032 N$6064 N$6063 "Straight Waveguide" sch_x=-99 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3033 N$6066 N$6065 "Straight Waveguide" sch_x=-99 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3034 N$6068 N$6067 "Straight Waveguide" sch_x=-99 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3035 N$6070 N$6069 "Straight Waveguide" sch_x=-99 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3036 N$6072 N$6071 "Straight Waveguide" sch_x=-99 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3037 N$6074 N$6073 "Straight Waveguide" sch_x=-99 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3038 N$6076 N$6075 "Straight Waveguide" sch_x=-99 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3039 N$6078 N$6077 "Straight Waveguide" sch_x=-99 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3040 N$6080 N$6079 "Straight Waveguide" sch_x=-99 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3041 N$6082 N$6081 "Straight Waveguide" sch_x=-99 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3042 N$6084 N$6083 "Straight Waveguide" sch_x=-99 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3043 N$6086 N$6085 "Straight Waveguide" sch_x=-99 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3044 N$6088 N$6087 "Straight Waveguide" sch_x=-99 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3045 N$6090 N$6089 "Straight Waveguide" sch_x=-99 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3046 N$6092 N$6091 "Straight Waveguide" sch_x=-99 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3047 N$6094 N$6093 "Straight Waveguide" sch_x=-99 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3048 N$6096 N$6095 "Straight Waveguide" sch_x=-99 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3049 N$6098 N$6097 "Straight Waveguide" sch_x=-99 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3050 N$6100 N$6099 "Straight Waveguide" sch_x=-99 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3051 N$6102 N$6101 "Straight Waveguide" sch_x=-99 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3052 N$6104 N$6103 "Straight Waveguide" sch_x=-99 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3053 N$6106 N$6105 "Straight Waveguide" sch_x=-99 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3054 N$6108 N$6107 "Straight Waveguide" sch_x=-99 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3055 N$6110 N$6109 "Straight Waveguide" sch_x=-97 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3056 N$6112 N$6111 "Straight Waveguide" sch_x=-97 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3057 N$6114 N$6113 "Straight Waveguide" sch_x=-97 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3058 N$6116 N$6115 "Straight Waveguide" sch_x=-97 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3059 N$6118 N$6117 "Straight Waveguide" sch_x=-97 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3060 N$6120 N$6119 "Straight Waveguide" sch_x=-97 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3061 N$6122 N$6121 "Straight Waveguide" sch_x=-97 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3062 N$6124 N$6123 "Straight Waveguide" sch_x=-97 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3063 N$6126 N$6125 "Straight Waveguide" sch_x=-97 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3064 N$6128 N$6127 "Straight Waveguide" sch_x=-97 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3065 N$6130 N$6129 "Straight Waveguide" sch_x=-97 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3066 N$6132 N$6131 "Straight Waveguide" sch_x=-97 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3067 N$6134 N$6133 "Straight Waveguide" sch_x=-97 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3068 N$6136 N$6135 "Straight Waveguide" sch_x=-97 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3069 N$6138 N$6137 "Straight Waveguide" sch_x=-97 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3070 N$6140 N$6139 "Straight Waveguide" sch_x=-97 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3071 N$6142 N$6141 "Straight Waveguide" sch_x=-97 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3072 N$6144 N$6143 "Straight Waveguide" sch_x=-97 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3073 N$6146 N$6145 "Straight Waveguide" sch_x=-97 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3074 N$6148 N$6147 "Straight Waveguide" sch_x=-97 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3075 N$6150 N$6149 "Straight Waveguide" sch_x=-97 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3076 N$6152 N$6151 "Straight Waveguide" sch_x=-97 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3077 N$6154 N$6153 "Straight Waveguide" sch_x=-97 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3078 N$6156 N$6155 "Straight Waveguide" sch_x=-97 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3079 N$6158 N$6157 "Straight Waveguide" sch_x=-97 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3080 N$6160 N$6159 "Straight Waveguide" sch_x=-97 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3081 N$6162 N$6161 "Straight Waveguide" sch_x=-97 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3082 N$6164 N$6163 "Straight Waveguide" sch_x=-97 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3083 N$6166 N$6165 "Straight Waveguide" sch_x=-97 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3084 N$6168 N$6167 "Straight Waveguide" sch_x=-97 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3085 N$6170 N$6169 "Straight Waveguide" sch_x=-97 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3086 N$6172 N$6171 "Straight Waveguide" sch_x=-97 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3087 N$6174 N$6173 "Straight Waveguide" sch_x=-97 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3088 N$6176 N$6175 "Straight Waveguide" sch_x=-97 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3089 N$6178 N$6177 "Straight Waveguide" sch_x=-95 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3090 N$6180 N$6179 "Straight Waveguide" sch_x=-95 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3091 N$6182 N$6181 "Straight Waveguide" sch_x=-95 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3092 N$6184 N$6183 "Straight Waveguide" sch_x=-95 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3093 N$6186 N$6185 "Straight Waveguide" sch_x=-95 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3094 N$6188 N$6187 "Straight Waveguide" sch_x=-95 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3095 N$6190 N$6189 "Straight Waveguide" sch_x=-95 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3096 N$6192 N$6191 "Straight Waveguide" sch_x=-95 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3097 N$6194 N$6193 "Straight Waveguide" sch_x=-95 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3098 N$6196 N$6195 "Straight Waveguide" sch_x=-95 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3099 N$6198 N$6197 "Straight Waveguide" sch_x=-95 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3100 N$6200 N$6199 "Straight Waveguide" sch_x=-95 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3101 N$6202 N$6201 "Straight Waveguide" sch_x=-95 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3102 N$6204 N$6203 "Straight Waveguide" sch_x=-95 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3103 N$6206 N$6205 "Straight Waveguide" sch_x=-95 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3104 N$6208 N$6207 "Straight Waveguide" sch_x=-95 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3105 N$6210 N$6209 "Straight Waveguide" sch_x=-95 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3106 N$6212 N$6211 "Straight Waveguide" sch_x=-95 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3107 N$6214 N$6213 "Straight Waveguide" sch_x=-95 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3108 N$6216 N$6215 "Straight Waveguide" sch_x=-95 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3109 N$6218 N$6217 "Straight Waveguide" sch_x=-95 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3110 N$6220 N$6219 "Straight Waveguide" sch_x=-95 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3111 N$6222 N$6221 "Straight Waveguide" sch_x=-95 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3112 N$6224 N$6223 "Straight Waveguide" sch_x=-95 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3113 N$6226 N$6225 "Straight Waveguide" sch_x=-95 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3114 N$6228 N$6227 "Straight Waveguide" sch_x=-95 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3115 N$6230 N$6229 "Straight Waveguide" sch_x=-95 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3116 N$6232 N$6231 "Straight Waveguide" sch_x=-95 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3117 N$6234 N$6233 "Straight Waveguide" sch_x=-95 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3118 N$6236 N$6235 "Straight Waveguide" sch_x=-95 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3119 N$6238 N$6237 "Straight Waveguide" sch_x=-95 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3120 N$6240 N$6239 "Straight Waveguide" sch_x=-95 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3121 N$6242 N$6241 "Straight Waveguide" sch_x=-93 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3122 N$6244 N$6243 "Straight Waveguide" sch_x=-93 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3123 N$6246 N$6245 "Straight Waveguide" sch_x=-93 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3124 N$6248 N$6247 "Straight Waveguide" sch_x=-93 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3125 N$6250 N$6249 "Straight Waveguide" sch_x=-93 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3126 N$6252 N$6251 "Straight Waveguide" sch_x=-93 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3127 N$6254 N$6253 "Straight Waveguide" sch_x=-93 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3128 N$6256 N$6255 "Straight Waveguide" sch_x=-93 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3129 N$6258 N$6257 "Straight Waveguide" sch_x=-93 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3130 N$6260 N$6259 "Straight Waveguide" sch_x=-93 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3131 N$6262 N$6261 "Straight Waveguide" sch_x=-93 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3132 N$6264 N$6263 "Straight Waveguide" sch_x=-93 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3133 N$6266 N$6265 "Straight Waveguide" sch_x=-93 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3134 N$6268 N$6267 "Straight Waveguide" sch_x=-93 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3135 N$6270 N$6269 "Straight Waveguide" sch_x=-93 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3136 N$6272 N$6271 "Straight Waveguide" sch_x=-93 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3137 N$6274 N$6273 "Straight Waveguide" sch_x=-93 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3138 N$6276 N$6275 "Straight Waveguide" sch_x=-93 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3139 N$6278 N$6277 "Straight Waveguide" sch_x=-93 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3140 N$6280 N$6279 "Straight Waveguide" sch_x=-93 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3141 N$6282 N$6281 "Straight Waveguide" sch_x=-93 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3142 N$6284 N$6283 "Straight Waveguide" sch_x=-93 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3143 N$6286 N$6285 "Straight Waveguide" sch_x=-93 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3144 N$6288 N$6287 "Straight Waveguide" sch_x=-93 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3145 N$6290 N$6289 "Straight Waveguide" sch_x=-93 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3146 N$6292 N$6291 "Straight Waveguide" sch_x=-93 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3147 N$6294 N$6293 "Straight Waveguide" sch_x=-93 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3148 N$6296 N$6295 "Straight Waveguide" sch_x=-93 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3149 N$6298 N$6297 "Straight Waveguide" sch_x=-93 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3150 N$6300 N$6299 "Straight Waveguide" sch_x=-93 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3151 N$6302 N$6301 "Straight Waveguide" sch_x=-91 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3152 N$6304 N$6303 "Straight Waveguide" sch_x=-91 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3153 N$6306 N$6305 "Straight Waveguide" sch_x=-91 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3154 N$6308 N$6307 "Straight Waveguide" sch_x=-91 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3155 N$6310 N$6309 "Straight Waveguide" sch_x=-91 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3156 N$6312 N$6311 "Straight Waveguide" sch_x=-91 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3157 N$6314 N$6313 "Straight Waveguide" sch_x=-91 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3158 N$6316 N$6315 "Straight Waveguide" sch_x=-91 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3159 N$6318 N$6317 "Straight Waveguide" sch_x=-91 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3160 N$6320 N$6319 "Straight Waveguide" sch_x=-91 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3161 N$6322 N$6321 "Straight Waveguide" sch_x=-91 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3162 N$6324 N$6323 "Straight Waveguide" sch_x=-91 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3163 N$6326 N$6325 "Straight Waveguide" sch_x=-91 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3164 N$6328 N$6327 "Straight Waveguide" sch_x=-91 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3165 N$6330 N$6329 "Straight Waveguide" sch_x=-91 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3166 N$6332 N$6331 "Straight Waveguide" sch_x=-91 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3167 N$6334 N$6333 "Straight Waveguide" sch_x=-91 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3168 N$6336 N$6335 "Straight Waveguide" sch_x=-91 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3169 N$6338 N$6337 "Straight Waveguide" sch_x=-91 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3170 N$6340 N$6339 "Straight Waveguide" sch_x=-91 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3171 N$6342 N$6341 "Straight Waveguide" sch_x=-91 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3172 N$6344 N$6343 "Straight Waveguide" sch_x=-91 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3173 N$6346 N$6345 "Straight Waveguide" sch_x=-91 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3174 N$6348 N$6347 "Straight Waveguide" sch_x=-91 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3175 N$6350 N$6349 "Straight Waveguide" sch_x=-91 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3176 N$6352 N$6351 "Straight Waveguide" sch_x=-91 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3177 N$6354 N$6353 "Straight Waveguide" sch_x=-91 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3178 N$6356 N$6355 "Straight Waveguide" sch_x=-91 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3179 N$6358 N$6357 "Straight Waveguide" sch_x=-89 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3180 N$6360 N$6359 "Straight Waveguide" sch_x=-89 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3181 N$6362 N$6361 "Straight Waveguide" sch_x=-89 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3182 N$6364 N$6363 "Straight Waveguide" sch_x=-89 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3183 N$6366 N$6365 "Straight Waveguide" sch_x=-89 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3184 N$6368 N$6367 "Straight Waveguide" sch_x=-89 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3185 N$6370 N$6369 "Straight Waveguide" sch_x=-89 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3186 N$6372 N$6371 "Straight Waveguide" sch_x=-89 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3187 N$6374 N$6373 "Straight Waveguide" sch_x=-89 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3188 N$6376 N$6375 "Straight Waveguide" sch_x=-89 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3189 N$6378 N$6377 "Straight Waveguide" sch_x=-89 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3190 N$6380 N$6379 "Straight Waveguide" sch_x=-89 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3191 N$6382 N$6381 "Straight Waveguide" sch_x=-89 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3192 N$6384 N$6383 "Straight Waveguide" sch_x=-89 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3193 N$6386 N$6385 "Straight Waveguide" sch_x=-89 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3194 N$6388 N$6387 "Straight Waveguide" sch_x=-89 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3195 N$6390 N$6389 "Straight Waveguide" sch_x=-89 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3196 N$6392 N$6391 "Straight Waveguide" sch_x=-89 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3197 N$6394 N$6393 "Straight Waveguide" sch_x=-89 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3198 N$6396 N$6395 "Straight Waveguide" sch_x=-89 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3199 N$6398 N$6397 "Straight Waveguide" sch_x=-89 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3200 N$6400 N$6399 "Straight Waveguide" sch_x=-89 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3201 N$6402 N$6401 "Straight Waveguide" sch_x=-89 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3202 N$6404 N$6403 "Straight Waveguide" sch_x=-89 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3203 N$6406 N$6405 "Straight Waveguide" sch_x=-89 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3204 N$6408 N$6407 "Straight Waveguide" sch_x=-89 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3205 N$6410 N$6409 "Straight Waveguide" sch_x=-87 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3206 N$6412 N$6411 "Straight Waveguide" sch_x=-87 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3207 N$6414 N$6413 "Straight Waveguide" sch_x=-87 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3208 N$6416 N$6415 "Straight Waveguide" sch_x=-87 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3209 N$6418 N$6417 "Straight Waveguide" sch_x=-87 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3210 N$6420 N$6419 "Straight Waveguide" sch_x=-87 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3211 N$6422 N$6421 "Straight Waveguide" sch_x=-87 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3212 N$6424 N$6423 "Straight Waveguide" sch_x=-87 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3213 N$6426 N$6425 "Straight Waveguide" sch_x=-87 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3214 N$6428 N$6427 "Straight Waveguide" sch_x=-87 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3215 N$6430 N$6429 "Straight Waveguide" sch_x=-87 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3216 N$6432 N$6431 "Straight Waveguide" sch_x=-87 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3217 N$6434 N$6433 "Straight Waveguide" sch_x=-87 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3218 N$6436 N$6435 "Straight Waveguide" sch_x=-87 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3219 N$6438 N$6437 "Straight Waveguide" sch_x=-87 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3220 N$6440 N$6439 "Straight Waveguide" sch_x=-87 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3221 N$6442 N$6441 "Straight Waveguide" sch_x=-87 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3222 N$6444 N$6443 "Straight Waveguide" sch_x=-87 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3223 N$6446 N$6445 "Straight Waveguide" sch_x=-87 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3224 N$6448 N$6447 "Straight Waveguide" sch_x=-87 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3225 N$6450 N$6449 "Straight Waveguide" sch_x=-87 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3226 N$6452 N$6451 "Straight Waveguide" sch_x=-87 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3227 N$6454 N$6453 "Straight Waveguide" sch_x=-87 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3228 N$6456 N$6455 "Straight Waveguide" sch_x=-87 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3229 N$6458 N$6457 "Straight Waveguide" sch_x=-85 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3230 N$6460 N$6459 "Straight Waveguide" sch_x=-85 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3231 N$6462 N$6461 "Straight Waveguide" sch_x=-85 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3232 N$6464 N$6463 "Straight Waveguide" sch_x=-85 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3233 N$6466 N$6465 "Straight Waveguide" sch_x=-85 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3234 N$6468 N$6467 "Straight Waveguide" sch_x=-85 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3235 N$6470 N$6469 "Straight Waveguide" sch_x=-85 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3236 N$6472 N$6471 "Straight Waveguide" sch_x=-85 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3237 N$6474 N$6473 "Straight Waveguide" sch_x=-85 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3238 N$6476 N$6475 "Straight Waveguide" sch_x=-85 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3239 N$6478 N$6477 "Straight Waveguide" sch_x=-85 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3240 N$6480 N$6479 "Straight Waveguide" sch_x=-85 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3241 N$6482 N$6481 "Straight Waveguide" sch_x=-85 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3242 N$6484 N$6483 "Straight Waveguide" sch_x=-85 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3243 N$6486 N$6485 "Straight Waveguide" sch_x=-85 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3244 N$6488 N$6487 "Straight Waveguide" sch_x=-85 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3245 N$6490 N$6489 "Straight Waveguide" sch_x=-85 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3246 N$6492 N$6491 "Straight Waveguide" sch_x=-85 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3247 N$6494 N$6493 "Straight Waveguide" sch_x=-85 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3248 N$6496 N$6495 "Straight Waveguide" sch_x=-85 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3249 N$6498 N$6497 "Straight Waveguide" sch_x=-85 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3250 N$6500 N$6499 "Straight Waveguide" sch_x=-85 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3251 N$6502 N$6501 "Straight Waveguide" sch_x=-83 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3252 N$6504 N$6503 "Straight Waveguide" sch_x=-83 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3253 N$6506 N$6505 "Straight Waveguide" sch_x=-83 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3254 N$6508 N$6507 "Straight Waveguide" sch_x=-83 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3255 N$6510 N$6509 "Straight Waveguide" sch_x=-83 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3256 N$6512 N$6511 "Straight Waveguide" sch_x=-83 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3257 N$6514 N$6513 "Straight Waveguide" sch_x=-83 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3258 N$6516 N$6515 "Straight Waveguide" sch_x=-83 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3259 N$6518 N$6517 "Straight Waveguide" sch_x=-83 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3260 N$6520 N$6519 "Straight Waveguide" sch_x=-83 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3261 N$6522 N$6521 "Straight Waveguide" sch_x=-83 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3262 N$6524 N$6523 "Straight Waveguide" sch_x=-83 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3263 N$6526 N$6525 "Straight Waveguide" sch_x=-83 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3264 N$6528 N$6527 "Straight Waveguide" sch_x=-83 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3265 N$6530 N$6529 "Straight Waveguide" sch_x=-83 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3266 N$6532 N$6531 "Straight Waveguide" sch_x=-83 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3267 N$6534 N$6533 "Straight Waveguide" sch_x=-83 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3268 N$6536 N$6535 "Straight Waveguide" sch_x=-83 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3269 N$6538 N$6537 "Straight Waveguide" sch_x=-83 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3270 N$6540 N$6539 "Straight Waveguide" sch_x=-83 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3271 N$6542 N$6541 "Straight Waveguide" sch_x=-81 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3272 N$6544 N$6543 "Straight Waveguide" sch_x=-81 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3273 N$6546 N$6545 "Straight Waveguide" sch_x=-81 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3274 N$6548 N$6547 "Straight Waveguide" sch_x=-81 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3275 N$6550 N$6549 "Straight Waveguide" sch_x=-81 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3276 N$6552 N$6551 "Straight Waveguide" sch_x=-81 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3277 N$6554 N$6553 "Straight Waveguide" sch_x=-81 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3278 N$6556 N$6555 "Straight Waveguide" sch_x=-81 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3279 N$6558 N$6557 "Straight Waveguide" sch_x=-81 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3280 N$6560 N$6559 "Straight Waveguide" sch_x=-81 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3281 N$6562 N$6561 "Straight Waveguide" sch_x=-81 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3282 N$6564 N$6563 "Straight Waveguide" sch_x=-81 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3283 N$6566 N$6565 "Straight Waveguide" sch_x=-81 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3284 N$6568 N$6567 "Straight Waveguide" sch_x=-81 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3285 N$6570 N$6569 "Straight Waveguide" sch_x=-81 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3286 N$6572 N$6571 "Straight Waveguide" sch_x=-81 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3287 N$6574 N$6573 "Straight Waveguide" sch_x=-81 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3288 N$6576 N$6575 "Straight Waveguide" sch_x=-81 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3289 N$6578 N$6577 "Straight Waveguide" sch_x=-79 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3290 N$6580 N$6579 "Straight Waveguide" sch_x=-79 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3291 N$6582 N$6581 "Straight Waveguide" sch_x=-79 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3292 N$6584 N$6583 "Straight Waveguide" sch_x=-79 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3293 N$6586 N$6585 "Straight Waveguide" sch_x=-79 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3294 N$6588 N$6587 "Straight Waveguide" sch_x=-79 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3295 N$6590 N$6589 "Straight Waveguide" sch_x=-79 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3296 N$6592 N$6591 "Straight Waveguide" sch_x=-79 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3297 N$6594 N$6593 "Straight Waveguide" sch_x=-79 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3298 N$6596 N$6595 "Straight Waveguide" sch_x=-79 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3299 N$6598 N$6597 "Straight Waveguide" sch_x=-79 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3300 N$6600 N$6599 "Straight Waveguide" sch_x=-79 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3301 N$6602 N$6601 "Straight Waveguide" sch_x=-79 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3302 N$6604 N$6603 "Straight Waveguide" sch_x=-79 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3303 N$6606 N$6605 "Straight Waveguide" sch_x=-79 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3304 N$6608 N$6607 "Straight Waveguide" sch_x=-79 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3305 N$6610 N$6609 "Straight Waveguide" sch_x=-77 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3306 N$6612 N$6611 "Straight Waveguide" sch_x=-77 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3307 N$6614 N$6613 "Straight Waveguide" sch_x=-77 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3308 N$6616 N$6615 "Straight Waveguide" sch_x=-77 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3309 N$6618 N$6617 "Straight Waveguide" sch_x=-77 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3310 N$6620 N$6619 "Straight Waveguide" sch_x=-77 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3311 N$6622 N$6621 "Straight Waveguide" sch_x=-77 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3312 N$6624 N$6623 "Straight Waveguide" sch_x=-77 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3313 N$6626 N$6625 "Straight Waveguide" sch_x=-77 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3314 N$6628 N$6627 "Straight Waveguide" sch_x=-77 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3315 N$6630 N$6629 "Straight Waveguide" sch_x=-77 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3316 N$6632 N$6631 "Straight Waveguide" sch_x=-77 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3317 N$6634 N$6633 "Straight Waveguide" sch_x=-77 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3318 N$6636 N$6635 "Straight Waveguide" sch_x=-77 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3319 N$6638 N$6637 "Straight Waveguide" sch_x=-75 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3320 N$6640 N$6639 "Straight Waveguide" sch_x=-75 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3321 N$6642 N$6641 "Straight Waveguide" sch_x=-75 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3322 N$6644 N$6643 "Straight Waveguide" sch_x=-75 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3323 N$6646 N$6645 "Straight Waveguide" sch_x=-75 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3324 N$6648 N$6647 "Straight Waveguide" sch_x=-75 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3325 N$6650 N$6649 "Straight Waveguide" sch_x=-75 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3326 N$6652 N$6651 "Straight Waveguide" sch_x=-75 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3327 N$6654 N$6653 "Straight Waveguide" sch_x=-75 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3328 N$6656 N$6655 "Straight Waveguide" sch_x=-75 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3329 N$6658 N$6657 "Straight Waveguide" sch_x=-75 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3330 N$6660 N$6659 "Straight Waveguide" sch_x=-75 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3331 N$6662 N$6661 "Straight Waveguide" sch_x=-73 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3332 N$6664 N$6663 "Straight Waveguide" sch_x=-73 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3333 N$6666 N$6665 "Straight Waveguide" sch_x=-73 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3334 N$6668 N$6667 "Straight Waveguide" sch_x=-73 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3335 N$6670 N$6669 "Straight Waveguide" sch_x=-73 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3336 N$6672 N$6671 "Straight Waveguide" sch_x=-73 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3337 N$6674 N$6673 "Straight Waveguide" sch_x=-73 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3338 N$6676 N$6675 "Straight Waveguide" sch_x=-73 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3339 N$6678 N$6677 "Straight Waveguide" sch_x=-73 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3340 N$6680 N$6679 "Straight Waveguide" sch_x=-73 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3341 N$6682 N$6681 "Straight Waveguide" sch_x=-71 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3342 N$6684 N$6683 "Straight Waveguide" sch_x=-71 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3343 N$6686 N$6685 "Straight Waveguide" sch_x=-71 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3344 N$6688 N$6687 "Straight Waveguide" sch_x=-71 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3345 N$6690 N$6689 "Straight Waveguide" sch_x=-71 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3346 N$6692 N$6691 "Straight Waveguide" sch_x=-71 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3347 N$6694 N$6693 "Straight Waveguide" sch_x=-71 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3348 N$6696 N$6695 "Straight Waveguide" sch_x=-71 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3349 N$6698 N$6697 "Straight Waveguide" sch_x=-69 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3350 N$6700 N$6699 "Straight Waveguide" sch_x=-69 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3351 N$6702 N$6701 "Straight Waveguide" sch_x=-69 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3352 N$6704 N$6703 "Straight Waveguide" sch_x=-69 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3353 N$6706 N$6705 "Straight Waveguide" sch_x=-69 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3354 N$6708 N$6707 "Straight Waveguide" sch_x=-69 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3355 N$6710 N$6709 "Straight Waveguide" sch_x=-67 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3356 N$6712 N$6711 "Straight Waveguide" sch_x=-67 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3357 N$6714 N$6713 "Straight Waveguide" sch_x=-67 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3358 N$6716 N$6715 "Straight Waveguide" sch_x=-67 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3359 N$6718 N$6717 "Straight Waveguide" sch_x=-65 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3360 N$6720 N$6719 "Straight Waveguide" sch_x=-65 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3361 N$6721 N$6722 "Straight Waveguide" sch_x=-93 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3362 N$6723 N$6724 "Straight Waveguide" sch_x=-92 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3363 N$6725 N$6726 "Straight Waveguide" sch_x=-91 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3364 N$6727 N$6728 "Straight Waveguide" sch_x=-90 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3365 N$6729 N$6730 "Straight Waveguide" sch_x=-89 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3366 N$6731 N$6732 "Straight Waveguide" sch_x=-88 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3367 N$6733 N$6734 "Straight Waveguide" sch_x=-87 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3368 N$6735 N$6736 "Straight Waveguide" sch_x=-86 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3369 N$6737 N$6738 "Straight Waveguide" sch_x=-85 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3370 N$6739 N$6740 "Straight Waveguide" sch_x=-84 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3371 N$6741 N$6742 "Straight Waveguide" sch_x=-83 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3372 N$6743 N$6744 "Straight Waveguide" sch_x=-82 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3373 N$6745 N$6746 "Straight Waveguide" sch_x=-81 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3374 N$6747 N$6748 "Straight Waveguide" sch_x=-80 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3375 N$6749 N$6750 "Straight Waveguide" sch_x=-79 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3376 N$6751 N$6752 "Straight Waveguide" sch_x=-78 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3377 N$6753 N$6754 "Straight Waveguide" sch_x=-77 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3378 N$6755 N$6756 "Straight Waveguide" sch_x=-76 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3379 N$6757 N$6758 "Straight Waveguide" sch_x=-75 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3380 N$6759 N$6760 "Straight Waveguide" sch_x=-74 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3381 N$6761 N$6762 "Straight Waveguide" sch_x=-73 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3382 N$6763 N$6764 "Straight Waveguide" sch_x=-72 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3383 N$6765 N$6766 "Straight Waveguide" sch_x=-71 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3384 N$6767 N$6768 "Straight Waveguide" sch_x=-70 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3385 N$6769 N$6770 "Straight Waveguide" sch_x=-69 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3386 N$6771 N$6772 "Straight Waveguide" sch_x=-68 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3387 N$6773 N$6774 "Straight Waveguide" sch_x=-67 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3388 N$6775 N$6776 "Straight Waveguide" sch_x=-66 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3389 N$6777 N$6778 "Straight Waveguide" sch_x=-65 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3390 N$6779 N$6780 "Straight Waveguide" sch_x=-64 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3391 N$6781 N$6782 "Straight Waveguide" sch_x=-63 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3392 N$6783 N$6784 "Straight Waveguide" sch_x=-63 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3393 N$6785 N$6786 "Straight Waveguide" sch_x=-64 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3394 N$6787 N$6788 "Straight Waveguide" sch_x=-65 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3395 N$6789 N$6790 "Straight Waveguide" sch_x=-66 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3396 N$6791 N$6792 "Straight Waveguide" sch_x=-67 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3397 N$6793 N$6794 "Straight Waveguide" sch_x=-68 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3398 N$6795 N$6796 "Straight Waveguide" sch_x=-69 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3399 N$6797 N$6798 "Straight Waveguide" sch_x=-70 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3400 N$6799 N$6800 "Straight Waveguide" sch_x=-71 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3401 N$6801 N$6802 "Straight Waveguide" sch_x=-72 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3402 N$6803 N$6804 "Straight Waveguide" sch_x=-73 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3403 N$6805 N$6806 "Straight Waveguide" sch_x=-74 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3404 N$6807 N$6808 "Straight Waveguide" sch_x=-75 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3405 N$6809 N$6810 "Straight Waveguide" sch_x=-76 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3406 N$6811 N$6812 "Straight Waveguide" sch_x=-77 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3407 N$6813 N$6814 "Straight Waveguide" sch_x=-78 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3408 N$6815 N$6816 "Straight Waveguide" sch_x=-79 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3409 N$6817 N$6818 "Straight Waveguide" sch_x=-80 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3410 N$6819 N$6820 "Straight Waveguide" sch_x=-81 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3411 N$6821 N$6822 "Straight Waveguide" sch_x=-82 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3412 N$6823 N$6824 "Straight Waveguide" sch_x=-83 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3413 N$6825 N$6826 "Straight Waveguide" sch_x=-84 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3414 N$6827 N$6828 "Straight Waveguide" sch_x=-85 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3415 N$6829 N$6830 "Straight Waveguide" sch_x=-86 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3416 N$6831 N$6832 "Straight Waveguide" sch_x=-87 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3417 N$6833 N$6834 "Straight Waveguide" sch_x=-88 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3418 N$6835 N$6836 "Straight Waveguide" sch_x=-89 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3419 N$6837 N$6838 "Straight Waveguide" sch_x=-90 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3420 N$6839 N$6840 "Straight Waveguide" sch_x=-91 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3421 N$6841 N$6842 "Straight Waveguide" sch_x=-92 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3422 N$6843 N$6844 "Straight Waveguide" sch_x=-93 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3423 N$6845 N$6846 "Straight Waveguide" sch_x=-94 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3424 N$6847 N$6848 "Straight Waveguide" sch_x=-94 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3425 N$6849 N$6850 "Straight Waveguide" sch_x=125 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3426 N$6851 N$6852 "Straight Waveguide" sch_x=125 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3427 N$6853 N$6854 "Straight Waveguide" sch_x=125 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3428 N$6855 N$6856 "Straight Waveguide" sch_x=125 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3429 N$6857 N$6858 "Straight Waveguide" sch_x=125 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3430 N$6859 N$6860 "Straight Waveguide" sch_x=125 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3431 N$6861 N$6862 "Straight Waveguide" sch_x=125 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3432 N$6863 N$6864 "Straight Waveguide" sch_x=125 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3433 N$6865 N$6866 "Straight Waveguide" sch_x=125 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3434 N$6867 N$6868 "Straight Waveguide" sch_x=125 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3435 N$6869 N$6870 "Straight Waveguide" sch_x=125 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3436 N$6871 N$6872 "Straight Waveguide" sch_x=125 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3437 N$6873 N$6874 "Straight Waveguide" sch_x=125 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3438 N$6875 N$6876 "Straight Waveguide" sch_x=125 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3439 N$6877 N$6878 "Straight Waveguide" sch_x=125 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3440 N$6879 N$6880 "Straight Waveguide" sch_x=125 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3441 N$6881 N$6882 "Straight Waveguide" sch_x=125 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3442 N$6883 N$6884 "Straight Waveguide" sch_x=125 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3443 N$6885 N$6886 "Straight Waveguide" sch_x=125 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3444 N$6887 N$6888 "Straight Waveguide" sch_x=125 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3445 N$6889 N$6890 "Straight Waveguide" sch_x=125 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3446 N$6891 N$6892 "Straight Waveguide" sch_x=125 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3447 N$6893 N$6894 "Straight Waveguide" sch_x=125 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3448 N$6895 N$6896 "Straight Waveguide" sch_x=125 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3449 N$6897 N$6898 "Straight Waveguide" sch_x=125 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3450 N$6899 N$6900 "Straight Waveguide" sch_x=125 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3451 N$6901 N$6902 "Straight Waveguide" sch_x=125 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3452 N$6903 N$6904 "Straight Waveguide" sch_x=125 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3453 N$6905 N$6906 "Straight Waveguide" sch_x=125 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3454 N$6907 N$6908 "Straight Waveguide" sch_x=125 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3455 N$6909 N$6910 "Straight Waveguide" sch_x=125 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3456 N$6911 N$6912 "Straight Waveguide" sch_x=125 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3457 N$6913 N$6914 "Straight Waveguide" sch_x=125 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3458 N$6915 N$6916 "Straight Waveguide" sch_x=125 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3459 N$6917 N$6918 "Straight Waveguide" sch_x=125 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3460 N$6919 N$6920 "Straight Waveguide" sch_x=125 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3461 N$6921 N$6922 "Straight Waveguide" sch_x=125 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3462 N$6923 N$6924 "Straight Waveguide" sch_x=125 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3463 N$6925 N$6926 "Straight Waveguide" sch_x=125 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3464 N$6927 N$6928 "Straight Waveguide" sch_x=125 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3465 N$6929 N$6930 "Straight Waveguide" sch_x=125 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3466 N$6931 N$6932 "Straight Waveguide" sch_x=125 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3467 N$6933 N$6934 "Straight Waveguide" sch_x=125 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3468 N$6935 N$6936 "Straight Waveguide" sch_x=125 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3469 N$6937 N$6938 "Straight Waveguide" sch_x=125 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3470 N$6939 N$6940 "Straight Waveguide" sch_x=125 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3471 N$6941 N$6942 "Straight Waveguide" sch_x=125 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3472 N$6943 N$6944 "Straight Waveguide" sch_x=125 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3473 N$6945 N$6946 "Straight Waveguide" sch_x=125 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3474 N$6947 N$6948 "Straight Waveguide" sch_x=125 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3475 N$6949 N$6950 "Straight Waveguide" sch_x=125 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3476 N$6951 N$6952 "Straight Waveguide" sch_x=125 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3477 N$6953 N$6954 "Straight Waveguide" sch_x=125 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3478 N$6955 N$6956 "Straight Waveguide" sch_x=125 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3479 N$6957 N$6958 "Straight Waveguide" sch_x=125 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3480 N$6959 N$6960 "Straight Waveguide" sch_x=125 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3481 N$6961 N$6962 "Straight Waveguide" sch_x=125 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3482 N$6963 N$6964 "Straight Waveguide" sch_x=125 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3483 N$6965 N$6966 "Straight Waveguide" sch_x=125 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3484 N$6967 N$6968 "Straight Waveguide" sch_x=125 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3485 N$6969 N$6970 "Straight Waveguide" sch_x=125 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3486 N$6971 N$6972 "Straight Waveguide" sch_x=125 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3487 N$6973 N$6974 "Straight Waveguide" sch_x=123 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3488 N$6975 N$6976 "Straight Waveguide" sch_x=123 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3489 N$6977 N$6978 "Straight Waveguide" sch_x=123 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3490 N$6979 N$6980 "Straight Waveguide" sch_x=123 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3491 N$6981 N$6982 "Straight Waveguide" sch_x=123 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3492 N$6983 N$6984 "Straight Waveguide" sch_x=123 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3493 N$6985 N$6986 "Straight Waveguide" sch_x=123 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3494 N$6987 N$6988 "Straight Waveguide" sch_x=123 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3495 N$6989 N$6990 "Straight Waveguide" sch_x=123 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3496 N$6991 N$6992 "Straight Waveguide" sch_x=123 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3497 N$6993 N$6994 "Straight Waveguide" sch_x=123 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3498 N$6995 N$6996 "Straight Waveguide" sch_x=123 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3499 N$6997 N$6998 "Straight Waveguide" sch_x=123 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3500 N$6999 N$7000 "Straight Waveguide" sch_x=123 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3501 N$7001 N$7002 "Straight Waveguide" sch_x=123 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3502 N$7003 N$7004 "Straight Waveguide" sch_x=123 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3503 N$7005 N$7006 "Straight Waveguide" sch_x=123 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3504 N$7007 N$7008 "Straight Waveguide" sch_x=123 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3505 N$7009 N$7010 "Straight Waveguide" sch_x=123 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3506 N$7011 N$7012 "Straight Waveguide" sch_x=123 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3507 N$7013 N$7014 "Straight Waveguide" sch_x=123 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3508 N$7015 N$7016 "Straight Waveguide" sch_x=123 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3509 N$7017 N$7018 "Straight Waveguide" sch_x=123 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3510 N$7019 N$7020 "Straight Waveguide" sch_x=123 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3511 N$7021 N$7022 "Straight Waveguide" sch_x=123 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3512 N$7023 N$7024 "Straight Waveguide" sch_x=123 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3513 N$7025 N$7026 "Straight Waveguide" sch_x=123 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3514 N$7027 N$7028 "Straight Waveguide" sch_x=123 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3515 N$7029 N$7030 "Straight Waveguide" sch_x=123 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3516 N$7031 N$7032 "Straight Waveguide" sch_x=123 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3517 N$7033 N$7034 "Straight Waveguide" sch_x=123 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3518 N$7035 N$7036 "Straight Waveguide" sch_x=123 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3519 N$7037 N$7038 "Straight Waveguide" sch_x=123 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3520 N$7039 N$7040 "Straight Waveguide" sch_x=123 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3521 N$7041 N$7042 "Straight Waveguide" sch_x=123 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3522 N$7043 N$7044 "Straight Waveguide" sch_x=123 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3523 N$7045 N$7046 "Straight Waveguide" sch_x=123 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3524 N$7047 N$7048 "Straight Waveguide" sch_x=123 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3525 N$7049 N$7050 "Straight Waveguide" sch_x=123 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3526 N$7051 N$7052 "Straight Waveguide" sch_x=123 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3527 N$7053 N$7054 "Straight Waveguide" sch_x=123 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3528 N$7055 N$7056 "Straight Waveguide" sch_x=123 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3529 N$7057 N$7058 "Straight Waveguide" sch_x=123 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3530 N$7059 N$7060 "Straight Waveguide" sch_x=123 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3531 N$7061 N$7062 "Straight Waveguide" sch_x=123 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3532 N$7063 N$7064 "Straight Waveguide" sch_x=123 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3533 N$7065 N$7066 "Straight Waveguide" sch_x=123 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3534 N$7067 N$7068 "Straight Waveguide" sch_x=123 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3535 N$7069 N$7070 "Straight Waveguide" sch_x=123 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3536 N$7071 N$7072 "Straight Waveguide" sch_x=123 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3537 N$7073 N$7074 "Straight Waveguide" sch_x=123 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3538 N$7075 N$7076 "Straight Waveguide" sch_x=123 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3539 N$7077 N$7078 "Straight Waveguide" sch_x=123 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3540 N$7079 N$7080 "Straight Waveguide" sch_x=123 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3541 N$7081 N$7082 "Straight Waveguide" sch_x=123 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3542 N$7083 N$7084 "Straight Waveguide" sch_x=123 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3543 N$7085 N$7086 "Straight Waveguide" sch_x=123 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3544 N$7087 N$7088 "Straight Waveguide" sch_x=123 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3545 N$7089 N$7090 "Straight Waveguide" sch_x=123 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3546 N$7091 N$7092 "Straight Waveguide" sch_x=123 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3547 N$7093 N$7094 "Straight Waveguide" sch_x=121 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3548 N$7095 N$7096 "Straight Waveguide" sch_x=121 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3549 N$7097 N$7098 "Straight Waveguide" sch_x=121 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3550 N$7099 N$7100 "Straight Waveguide" sch_x=121 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3551 N$7101 N$7102 "Straight Waveguide" sch_x=121 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3552 N$7103 N$7104 "Straight Waveguide" sch_x=121 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3553 N$7105 N$7106 "Straight Waveguide" sch_x=121 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3554 N$7107 N$7108 "Straight Waveguide" sch_x=121 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3555 N$7109 N$7110 "Straight Waveguide" sch_x=121 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3556 N$7111 N$7112 "Straight Waveguide" sch_x=121 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3557 N$7113 N$7114 "Straight Waveguide" sch_x=121 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3558 N$7115 N$7116 "Straight Waveguide" sch_x=121 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3559 N$7117 N$7118 "Straight Waveguide" sch_x=121 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3560 N$7119 N$7120 "Straight Waveguide" sch_x=121 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3561 N$7121 N$7122 "Straight Waveguide" sch_x=121 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3562 N$7123 N$7124 "Straight Waveguide" sch_x=121 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3563 N$7125 N$7126 "Straight Waveguide" sch_x=121 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3564 N$7127 N$7128 "Straight Waveguide" sch_x=121 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3565 N$7129 N$7130 "Straight Waveguide" sch_x=121 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3566 N$7131 N$7132 "Straight Waveguide" sch_x=121 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3567 N$7133 N$7134 "Straight Waveguide" sch_x=121 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3568 N$7135 N$7136 "Straight Waveguide" sch_x=121 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3569 N$7137 N$7138 "Straight Waveguide" sch_x=121 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3570 N$7139 N$7140 "Straight Waveguide" sch_x=121 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3571 N$7141 N$7142 "Straight Waveguide" sch_x=121 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3572 N$7143 N$7144 "Straight Waveguide" sch_x=121 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3573 N$7145 N$7146 "Straight Waveguide" sch_x=121 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3574 N$7147 N$7148 "Straight Waveguide" sch_x=121 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3575 N$7149 N$7150 "Straight Waveguide" sch_x=121 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3576 N$7151 N$7152 "Straight Waveguide" sch_x=121 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3577 N$7153 N$7154 "Straight Waveguide" sch_x=121 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3578 N$7155 N$7156 "Straight Waveguide" sch_x=121 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3579 N$7157 N$7158 "Straight Waveguide" sch_x=121 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3580 N$7159 N$7160 "Straight Waveguide" sch_x=121 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3581 N$7161 N$7162 "Straight Waveguide" sch_x=121 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3582 N$7163 N$7164 "Straight Waveguide" sch_x=121 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3583 N$7165 N$7166 "Straight Waveguide" sch_x=121 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3584 N$7167 N$7168 "Straight Waveguide" sch_x=121 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3585 N$7169 N$7170 "Straight Waveguide" sch_x=121 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3586 N$7171 N$7172 "Straight Waveguide" sch_x=121 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3587 N$7173 N$7174 "Straight Waveguide" sch_x=121 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3588 N$7175 N$7176 "Straight Waveguide" sch_x=121 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3589 N$7177 N$7178 "Straight Waveguide" sch_x=121 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3590 N$7179 N$7180 "Straight Waveguide" sch_x=121 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3591 N$7181 N$7182 "Straight Waveguide" sch_x=121 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3592 N$7183 N$7184 "Straight Waveguide" sch_x=121 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3593 N$7185 N$7186 "Straight Waveguide" sch_x=121 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3594 N$7187 N$7188 "Straight Waveguide" sch_x=121 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3595 N$7189 N$7190 "Straight Waveguide" sch_x=121 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3596 N$7191 N$7192 "Straight Waveguide" sch_x=121 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3597 N$7193 N$7194 "Straight Waveguide" sch_x=121 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3598 N$7195 N$7196 "Straight Waveguide" sch_x=121 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3599 N$7197 N$7198 "Straight Waveguide" sch_x=121 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3600 N$7199 N$7200 "Straight Waveguide" sch_x=121 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3601 N$7201 N$7202 "Straight Waveguide" sch_x=121 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3602 N$7203 N$7204 "Straight Waveguide" sch_x=121 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3603 N$7205 N$7206 "Straight Waveguide" sch_x=121 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3604 N$7207 N$7208 "Straight Waveguide" sch_x=121 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3605 N$7209 N$7210 "Straight Waveguide" sch_x=119 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3606 N$7211 N$7212 "Straight Waveguide" sch_x=119 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3607 N$7213 N$7214 "Straight Waveguide" sch_x=119 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3608 N$7215 N$7216 "Straight Waveguide" sch_x=119 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3609 N$7217 N$7218 "Straight Waveguide" sch_x=119 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3610 N$7219 N$7220 "Straight Waveguide" sch_x=119 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3611 N$7221 N$7222 "Straight Waveguide" sch_x=119 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3612 N$7223 N$7224 "Straight Waveguide" sch_x=119 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3613 N$7225 N$7226 "Straight Waveguide" sch_x=119 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3614 N$7227 N$7228 "Straight Waveguide" sch_x=119 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3615 N$7229 N$7230 "Straight Waveguide" sch_x=119 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3616 N$7231 N$7232 "Straight Waveguide" sch_x=119 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3617 N$7233 N$7234 "Straight Waveguide" sch_x=119 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3618 N$7235 N$7236 "Straight Waveguide" sch_x=119 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3619 N$7237 N$7238 "Straight Waveguide" sch_x=119 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3620 N$7239 N$7240 "Straight Waveguide" sch_x=119 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3621 N$7241 N$7242 "Straight Waveguide" sch_x=119 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3622 N$7243 N$7244 "Straight Waveguide" sch_x=119 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3623 N$7245 N$7246 "Straight Waveguide" sch_x=119 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3624 N$7247 N$7248 "Straight Waveguide" sch_x=119 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3625 N$7249 N$7250 "Straight Waveguide" sch_x=119 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3626 N$7251 N$7252 "Straight Waveguide" sch_x=119 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3627 N$7253 N$7254 "Straight Waveguide" sch_x=119 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3628 N$7255 N$7256 "Straight Waveguide" sch_x=119 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3629 N$7257 N$7258 "Straight Waveguide" sch_x=119 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3630 N$7259 N$7260 "Straight Waveguide" sch_x=119 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3631 N$7261 N$7262 "Straight Waveguide" sch_x=119 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3632 N$7263 N$7264 "Straight Waveguide" sch_x=119 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3633 N$7265 N$7266 "Straight Waveguide" sch_x=119 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3634 N$7267 N$7268 "Straight Waveguide" sch_x=119 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3635 N$7269 N$7270 "Straight Waveguide" sch_x=119 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3636 N$7271 N$7272 "Straight Waveguide" sch_x=119 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3637 N$7273 N$7274 "Straight Waveguide" sch_x=119 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3638 N$7275 N$7276 "Straight Waveguide" sch_x=119 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3639 N$7277 N$7278 "Straight Waveguide" sch_x=119 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3640 N$7279 N$7280 "Straight Waveguide" sch_x=119 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3641 N$7281 N$7282 "Straight Waveguide" sch_x=119 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3642 N$7283 N$7284 "Straight Waveguide" sch_x=119 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3643 N$7285 N$7286 "Straight Waveguide" sch_x=119 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3644 N$7287 N$7288 "Straight Waveguide" sch_x=119 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3645 N$7289 N$7290 "Straight Waveguide" sch_x=119 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3646 N$7291 N$7292 "Straight Waveguide" sch_x=119 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3647 N$7293 N$7294 "Straight Waveguide" sch_x=119 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3648 N$7295 N$7296 "Straight Waveguide" sch_x=119 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3649 N$7297 N$7298 "Straight Waveguide" sch_x=119 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3650 N$7299 N$7300 "Straight Waveguide" sch_x=119 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3651 N$7301 N$7302 "Straight Waveguide" sch_x=119 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3652 N$7303 N$7304 "Straight Waveguide" sch_x=119 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3653 N$7305 N$7306 "Straight Waveguide" sch_x=119 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3654 N$7307 N$7308 "Straight Waveguide" sch_x=119 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3655 N$7309 N$7310 "Straight Waveguide" sch_x=119 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3656 N$7311 N$7312 "Straight Waveguide" sch_x=119 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3657 N$7313 N$7314 "Straight Waveguide" sch_x=119 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3658 N$7315 N$7316 "Straight Waveguide" sch_x=119 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3659 N$7317 N$7318 "Straight Waveguide" sch_x=119 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3660 N$7319 N$7320 "Straight Waveguide" sch_x=119 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3661 N$7321 N$7322 "Straight Waveguide" sch_x=117 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3662 N$7323 N$7324 "Straight Waveguide" sch_x=117 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3663 N$7325 N$7326 "Straight Waveguide" sch_x=117 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3664 N$7327 N$7328 "Straight Waveguide" sch_x=117 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3665 N$7329 N$7330 "Straight Waveguide" sch_x=117 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3666 N$7331 N$7332 "Straight Waveguide" sch_x=117 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3667 N$7333 N$7334 "Straight Waveguide" sch_x=117 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3668 N$7335 N$7336 "Straight Waveguide" sch_x=117 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3669 N$7337 N$7338 "Straight Waveguide" sch_x=117 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3670 N$7339 N$7340 "Straight Waveguide" sch_x=117 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3671 N$7341 N$7342 "Straight Waveguide" sch_x=117 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3672 N$7343 N$7344 "Straight Waveguide" sch_x=117 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3673 N$7345 N$7346 "Straight Waveguide" sch_x=117 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3674 N$7347 N$7348 "Straight Waveguide" sch_x=117 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3675 N$7349 N$7350 "Straight Waveguide" sch_x=117 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3676 N$7351 N$7352 "Straight Waveguide" sch_x=117 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3677 N$7353 N$7354 "Straight Waveguide" sch_x=117 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3678 N$7355 N$7356 "Straight Waveguide" sch_x=117 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3679 N$7357 N$7358 "Straight Waveguide" sch_x=117 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3680 N$7359 N$7360 "Straight Waveguide" sch_x=117 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3681 N$7361 N$7362 "Straight Waveguide" sch_x=117 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3682 N$7363 N$7364 "Straight Waveguide" sch_x=117 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3683 N$7365 N$7366 "Straight Waveguide" sch_x=117 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3684 N$7367 N$7368 "Straight Waveguide" sch_x=117 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3685 N$7369 N$7370 "Straight Waveguide" sch_x=117 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3686 N$7371 N$7372 "Straight Waveguide" sch_x=117 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3687 N$7373 N$7374 "Straight Waveguide" sch_x=117 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3688 N$7375 N$7376 "Straight Waveguide" sch_x=117 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3689 N$7377 N$7378 "Straight Waveguide" sch_x=117 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3690 N$7379 N$7380 "Straight Waveguide" sch_x=117 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3691 N$7381 N$7382 "Straight Waveguide" sch_x=117 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3692 N$7383 N$7384 "Straight Waveguide" sch_x=117 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3693 N$7385 N$7386 "Straight Waveguide" sch_x=117 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3694 N$7387 N$7388 "Straight Waveguide" sch_x=117 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3695 N$7389 N$7390 "Straight Waveguide" sch_x=117 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3696 N$7391 N$7392 "Straight Waveguide" sch_x=117 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3697 N$7393 N$7394 "Straight Waveguide" sch_x=117 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3698 N$7395 N$7396 "Straight Waveguide" sch_x=117 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3699 N$7397 N$7398 "Straight Waveguide" sch_x=117 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3700 N$7399 N$7400 "Straight Waveguide" sch_x=117 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3701 N$7401 N$7402 "Straight Waveguide" sch_x=117 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3702 N$7403 N$7404 "Straight Waveguide" sch_x=117 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3703 N$7405 N$7406 "Straight Waveguide" sch_x=117 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3704 N$7407 N$7408 "Straight Waveguide" sch_x=117 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3705 N$7409 N$7410 "Straight Waveguide" sch_x=117 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3706 N$7411 N$7412 "Straight Waveguide" sch_x=117 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3707 N$7413 N$7414 "Straight Waveguide" sch_x=117 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3708 N$7415 N$7416 "Straight Waveguide" sch_x=117 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3709 N$7417 N$7418 "Straight Waveguide" sch_x=117 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3710 N$7419 N$7420 "Straight Waveguide" sch_x=117 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3711 N$7421 N$7422 "Straight Waveguide" sch_x=117 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3712 N$7423 N$7424 "Straight Waveguide" sch_x=117 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3713 N$7425 N$7426 "Straight Waveguide" sch_x=117 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3714 N$7427 N$7428 "Straight Waveguide" sch_x=117 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3715 N$7429 N$7430 "Straight Waveguide" sch_x=115 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3716 N$7431 N$7432 "Straight Waveguide" sch_x=115 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3717 N$7433 N$7434 "Straight Waveguide" sch_x=115 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3718 N$7435 N$7436 "Straight Waveguide" sch_x=115 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3719 N$7437 N$7438 "Straight Waveguide" sch_x=115 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3720 N$7439 N$7440 "Straight Waveguide" sch_x=115 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3721 N$7441 N$7442 "Straight Waveguide" sch_x=115 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3722 N$7443 N$7444 "Straight Waveguide" sch_x=115 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3723 N$7445 N$7446 "Straight Waveguide" sch_x=115 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3724 N$7447 N$7448 "Straight Waveguide" sch_x=115 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3725 N$7449 N$7450 "Straight Waveguide" sch_x=115 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3726 N$7451 N$7452 "Straight Waveguide" sch_x=115 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3727 N$7453 N$7454 "Straight Waveguide" sch_x=115 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3728 N$7455 N$7456 "Straight Waveguide" sch_x=115 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3729 N$7457 N$7458 "Straight Waveguide" sch_x=115 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3730 N$7459 N$7460 "Straight Waveguide" sch_x=115 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3731 N$7461 N$7462 "Straight Waveguide" sch_x=115 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3732 N$7463 N$7464 "Straight Waveguide" sch_x=115 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3733 N$7465 N$7466 "Straight Waveguide" sch_x=115 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3734 N$7467 N$7468 "Straight Waveguide" sch_x=115 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3735 N$7469 N$7470 "Straight Waveguide" sch_x=115 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3736 N$7471 N$7472 "Straight Waveguide" sch_x=115 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3737 N$7473 N$7474 "Straight Waveguide" sch_x=115 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3738 N$7475 N$7476 "Straight Waveguide" sch_x=115 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3739 N$7477 N$7478 "Straight Waveguide" sch_x=115 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3740 N$7479 N$7480 "Straight Waveguide" sch_x=115 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3741 N$7481 N$7482 "Straight Waveguide" sch_x=115 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3742 N$7483 N$7484 "Straight Waveguide" sch_x=115 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3743 N$7485 N$7486 "Straight Waveguide" sch_x=115 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3744 N$7487 N$7488 "Straight Waveguide" sch_x=115 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3745 N$7489 N$7490 "Straight Waveguide" sch_x=115 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3746 N$7491 N$7492 "Straight Waveguide" sch_x=115 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3747 N$7493 N$7494 "Straight Waveguide" sch_x=115 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3748 N$7495 N$7496 "Straight Waveguide" sch_x=115 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3749 N$7497 N$7498 "Straight Waveguide" sch_x=115 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3750 N$7499 N$7500 "Straight Waveguide" sch_x=115 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3751 N$7501 N$7502 "Straight Waveguide" sch_x=115 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3752 N$7503 N$7504 "Straight Waveguide" sch_x=115 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3753 N$7505 N$7506 "Straight Waveguide" sch_x=115 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3754 N$7507 N$7508 "Straight Waveguide" sch_x=115 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3755 N$7509 N$7510 "Straight Waveguide" sch_x=115 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3756 N$7511 N$7512 "Straight Waveguide" sch_x=115 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3757 N$7513 N$7514 "Straight Waveguide" sch_x=115 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3758 N$7515 N$7516 "Straight Waveguide" sch_x=115 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3759 N$7517 N$7518 "Straight Waveguide" sch_x=115 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3760 N$7519 N$7520 "Straight Waveguide" sch_x=115 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3761 N$7521 N$7522 "Straight Waveguide" sch_x=115 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3762 N$7523 N$7524 "Straight Waveguide" sch_x=115 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3763 N$7525 N$7526 "Straight Waveguide" sch_x=115 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3764 N$7527 N$7528 "Straight Waveguide" sch_x=115 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3765 N$7529 N$7530 "Straight Waveguide" sch_x=115 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3766 N$7531 N$7532 "Straight Waveguide" sch_x=115 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3767 N$7533 N$7534 "Straight Waveguide" sch_x=113 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3768 N$7535 N$7536 "Straight Waveguide" sch_x=113 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3769 N$7537 N$7538 "Straight Waveguide" sch_x=113 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3770 N$7539 N$7540 "Straight Waveguide" sch_x=113 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3771 N$7541 N$7542 "Straight Waveguide" sch_x=113 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3772 N$7543 N$7544 "Straight Waveguide" sch_x=113 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3773 N$7545 N$7546 "Straight Waveguide" sch_x=113 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3774 N$7547 N$7548 "Straight Waveguide" sch_x=113 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3775 N$7549 N$7550 "Straight Waveguide" sch_x=113 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3776 N$7551 N$7552 "Straight Waveguide" sch_x=113 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3777 N$7553 N$7554 "Straight Waveguide" sch_x=113 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3778 N$7555 N$7556 "Straight Waveguide" sch_x=113 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3779 N$7557 N$7558 "Straight Waveguide" sch_x=113 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3780 N$7559 N$7560 "Straight Waveguide" sch_x=113 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3781 N$7561 N$7562 "Straight Waveguide" sch_x=113 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3782 N$7563 N$7564 "Straight Waveguide" sch_x=113 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3783 N$7565 N$7566 "Straight Waveguide" sch_x=113 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3784 N$7567 N$7568 "Straight Waveguide" sch_x=113 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3785 N$7569 N$7570 "Straight Waveguide" sch_x=113 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3786 N$7571 N$7572 "Straight Waveguide" sch_x=113 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3787 N$7573 N$7574 "Straight Waveguide" sch_x=113 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3788 N$7575 N$7576 "Straight Waveguide" sch_x=113 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3789 N$7577 N$7578 "Straight Waveguide" sch_x=113 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3790 N$7579 N$7580 "Straight Waveguide" sch_x=113 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3791 N$7581 N$7582 "Straight Waveguide" sch_x=113 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3792 N$7583 N$7584 "Straight Waveguide" sch_x=113 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3793 N$7585 N$7586 "Straight Waveguide" sch_x=113 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3794 N$7587 N$7588 "Straight Waveguide" sch_x=113 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3795 N$7589 N$7590 "Straight Waveguide" sch_x=113 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3796 N$7591 N$7592 "Straight Waveguide" sch_x=113 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3797 N$7593 N$7594 "Straight Waveguide" sch_x=113 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3798 N$7595 N$7596 "Straight Waveguide" sch_x=113 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3799 N$7597 N$7598 "Straight Waveguide" sch_x=113 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3800 N$7599 N$7600 "Straight Waveguide" sch_x=113 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3801 N$7601 N$7602 "Straight Waveguide" sch_x=113 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3802 N$7603 N$7604 "Straight Waveguide" sch_x=113 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3803 N$7605 N$7606 "Straight Waveguide" sch_x=113 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3804 N$7607 N$7608 "Straight Waveguide" sch_x=113 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3805 N$7609 N$7610 "Straight Waveguide" sch_x=113 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3806 N$7611 N$7612 "Straight Waveguide" sch_x=113 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3807 N$7613 N$7614 "Straight Waveguide" sch_x=113 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3808 N$7615 N$7616 "Straight Waveguide" sch_x=113 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3809 N$7617 N$7618 "Straight Waveguide" sch_x=113 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3810 N$7619 N$7620 "Straight Waveguide" sch_x=113 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3811 N$7621 N$7622 "Straight Waveguide" sch_x=113 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3812 N$7623 N$7624 "Straight Waveguide" sch_x=113 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3813 N$7625 N$7626 "Straight Waveguide" sch_x=113 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3814 N$7627 N$7628 "Straight Waveguide" sch_x=113 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3815 N$7629 N$7630 "Straight Waveguide" sch_x=113 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3816 N$7631 N$7632 "Straight Waveguide" sch_x=113 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3817 N$7633 N$7634 "Straight Waveguide" sch_x=111 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3818 N$7635 N$7636 "Straight Waveguide" sch_x=111 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3819 N$7637 N$7638 "Straight Waveguide" sch_x=111 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3820 N$7639 N$7640 "Straight Waveguide" sch_x=111 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3821 N$7641 N$7642 "Straight Waveguide" sch_x=111 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3822 N$7643 N$7644 "Straight Waveguide" sch_x=111 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3823 N$7645 N$7646 "Straight Waveguide" sch_x=111 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3824 N$7647 N$7648 "Straight Waveguide" sch_x=111 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3825 N$7649 N$7650 "Straight Waveguide" sch_x=111 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3826 N$7651 N$7652 "Straight Waveguide" sch_x=111 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3827 N$7653 N$7654 "Straight Waveguide" sch_x=111 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3828 N$7655 N$7656 "Straight Waveguide" sch_x=111 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3829 N$7657 N$7658 "Straight Waveguide" sch_x=111 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3830 N$7659 N$7660 "Straight Waveguide" sch_x=111 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3831 N$7661 N$7662 "Straight Waveguide" sch_x=111 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3832 N$7663 N$7664 "Straight Waveguide" sch_x=111 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3833 N$7665 N$7666 "Straight Waveguide" sch_x=111 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3834 N$7667 N$7668 "Straight Waveguide" sch_x=111 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3835 N$7669 N$7670 "Straight Waveguide" sch_x=111 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3836 N$7671 N$7672 "Straight Waveguide" sch_x=111 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3837 N$7673 N$7674 "Straight Waveguide" sch_x=111 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3838 N$7675 N$7676 "Straight Waveguide" sch_x=111 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3839 N$7677 N$7678 "Straight Waveguide" sch_x=111 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3840 N$7679 N$7680 "Straight Waveguide" sch_x=111 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3841 N$7681 N$7682 "Straight Waveguide" sch_x=111 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3842 N$7683 N$7684 "Straight Waveguide" sch_x=111 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3843 N$7685 N$7686 "Straight Waveguide" sch_x=111 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3844 N$7687 N$7688 "Straight Waveguide" sch_x=111 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3845 N$7689 N$7690 "Straight Waveguide" sch_x=111 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3846 N$7691 N$7692 "Straight Waveguide" sch_x=111 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3847 N$7693 N$7694 "Straight Waveguide" sch_x=111 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3848 N$7695 N$7696 "Straight Waveguide" sch_x=111 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3849 N$7697 N$7698 "Straight Waveguide" sch_x=111 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3850 N$7699 N$7700 "Straight Waveguide" sch_x=111 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3851 N$7701 N$7702 "Straight Waveguide" sch_x=111 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3852 N$7703 N$7704 "Straight Waveguide" sch_x=111 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3853 N$7705 N$7706 "Straight Waveguide" sch_x=111 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3854 N$7707 N$7708 "Straight Waveguide" sch_x=111 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3855 N$7709 N$7710 "Straight Waveguide" sch_x=111 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3856 N$7711 N$7712 "Straight Waveguide" sch_x=111 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3857 N$7713 N$7714 "Straight Waveguide" sch_x=111 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3858 N$7715 N$7716 "Straight Waveguide" sch_x=111 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3859 N$7717 N$7718 "Straight Waveguide" sch_x=111 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3860 N$7719 N$7720 "Straight Waveguide" sch_x=111 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3861 N$7721 N$7722 "Straight Waveguide" sch_x=111 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3862 N$7723 N$7724 "Straight Waveguide" sch_x=111 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3863 N$7725 N$7726 "Straight Waveguide" sch_x=111 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3864 N$7727 N$7728 "Straight Waveguide" sch_x=111 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3865 N$7729 N$7730 "Straight Waveguide" sch_x=109 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3866 N$7731 N$7732 "Straight Waveguide" sch_x=109 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3867 N$7733 N$7734 "Straight Waveguide" sch_x=109 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3868 N$7735 N$7736 "Straight Waveguide" sch_x=109 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3869 N$7737 N$7738 "Straight Waveguide" sch_x=109 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3870 N$7739 N$7740 "Straight Waveguide" sch_x=109 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3871 N$7741 N$7742 "Straight Waveguide" sch_x=109 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3872 N$7743 N$7744 "Straight Waveguide" sch_x=109 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3873 N$7745 N$7746 "Straight Waveguide" sch_x=109 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3874 N$7747 N$7748 "Straight Waveguide" sch_x=109 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3875 N$7749 N$7750 "Straight Waveguide" sch_x=109 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3876 N$7751 N$7752 "Straight Waveguide" sch_x=109 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3877 N$7753 N$7754 "Straight Waveguide" sch_x=109 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3878 N$7755 N$7756 "Straight Waveguide" sch_x=109 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3879 N$7757 N$7758 "Straight Waveguide" sch_x=109 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3880 N$7759 N$7760 "Straight Waveguide" sch_x=109 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3881 N$7761 N$7762 "Straight Waveguide" sch_x=109 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3882 N$7763 N$7764 "Straight Waveguide" sch_x=109 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3883 N$7765 N$7766 "Straight Waveguide" sch_x=109 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3884 N$7767 N$7768 "Straight Waveguide" sch_x=109 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3885 N$7769 N$7770 "Straight Waveguide" sch_x=109 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3886 N$7771 N$7772 "Straight Waveguide" sch_x=109 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3887 N$7773 N$7774 "Straight Waveguide" sch_x=109 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3888 N$7775 N$7776 "Straight Waveguide" sch_x=109 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3889 N$7777 N$7778 "Straight Waveguide" sch_x=109 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3890 N$7779 N$7780 "Straight Waveguide" sch_x=109 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3891 N$7781 N$7782 "Straight Waveguide" sch_x=109 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3892 N$7783 N$7784 "Straight Waveguide" sch_x=109 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3893 N$7785 N$7786 "Straight Waveguide" sch_x=109 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3894 N$7787 N$7788 "Straight Waveguide" sch_x=109 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3895 N$7789 N$7790 "Straight Waveguide" sch_x=109 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3896 N$7791 N$7792 "Straight Waveguide" sch_x=109 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3897 N$7793 N$7794 "Straight Waveguide" sch_x=109 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3898 N$7795 N$7796 "Straight Waveguide" sch_x=109 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3899 N$7797 N$7798 "Straight Waveguide" sch_x=109 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3900 N$7799 N$7800 "Straight Waveguide" sch_x=109 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3901 N$7801 N$7802 "Straight Waveguide" sch_x=109 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3902 N$7803 N$7804 "Straight Waveguide" sch_x=109 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3903 N$7805 N$7806 "Straight Waveguide" sch_x=109 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3904 N$7807 N$7808 "Straight Waveguide" sch_x=109 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3905 N$7809 N$7810 "Straight Waveguide" sch_x=109 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3906 N$7811 N$7812 "Straight Waveguide" sch_x=109 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3907 N$7813 N$7814 "Straight Waveguide" sch_x=109 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3908 N$7815 N$7816 "Straight Waveguide" sch_x=109 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3909 N$7817 N$7818 "Straight Waveguide" sch_x=109 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3910 N$7819 N$7820 "Straight Waveguide" sch_x=109 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3911 N$7821 N$7822 "Straight Waveguide" sch_x=107 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3912 N$7823 N$7824 "Straight Waveguide" sch_x=107 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3913 N$7825 N$7826 "Straight Waveguide" sch_x=107 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3914 N$7827 N$7828 "Straight Waveguide" sch_x=107 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3915 N$7829 N$7830 "Straight Waveguide" sch_x=107 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3916 N$7831 N$7832 "Straight Waveguide" sch_x=107 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3917 N$7833 N$7834 "Straight Waveguide" sch_x=107 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3918 N$7835 N$7836 "Straight Waveguide" sch_x=107 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3919 N$7837 N$7838 "Straight Waveguide" sch_x=107 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3920 N$7839 N$7840 "Straight Waveguide" sch_x=107 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3921 N$7841 N$7842 "Straight Waveguide" sch_x=107 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3922 N$7843 N$7844 "Straight Waveguide" sch_x=107 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3923 N$7845 N$7846 "Straight Waveguide" sch_x=107 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3924 N$7847 N$7848 "Straight Waveguide" sch_x=107 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3925 N$7849 N$7850 "Straight Waveguide" sch_x=107 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3926 N$7851 N$7852 "Straight Waveguide" sch_x=107 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3927 N$7853 N$7854 "Straight Waveguide" sch_x=107 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3928 N$7855 N$7856 "Straight Waveguide" sch_x=107 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3929 N$7857 N$7858 "Straight Waveguide" sch_x=107 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3930 N$7859 N$7860 "Straight Waveguide" sch_x=107 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3931 N$7861 N$7862 "Straight Waveguide" sch_x=107 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3932 N$7863 N$7864 "Straight Waveguide" sch_x=107 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3933 N$7865 N$7866 "Straight Waveguide" sch_x=107 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3934 N$7867 N$7868 "Straight Waveguide" sch_x=107 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3935 N$7869 N$7870 "Straight Waveguide" sch_x=107 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3936 N$7871 N$7872 "Straight Waveguide" sch_x=107 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3937 N$7873 N$7874 "Straight Waveguide" sch_x=107 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3938 N$7875 N$7876 "Straight Waveguide" sch_x=107 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3939 N$7877 N$7878 "Straight Waveguide" sch_x=107 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3940 N$7879 N$7880 "Straight Waveguide" sch_x=107 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3941 N$7881 N$7882 "Straight Waveguide" sch_x=107 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3942 N$7883 N$7884 "Straight Waveguide" sch_x=107 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3943 N$7885 N$7886 "Straight Waveguide" sch_x=107 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3944 N$7887 N$7888 "Straight Waveguide" sch_x=107 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3945 N$7889 N$7890 "Straight Waveguide" sch_x=107 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3946 N$7891 N$7892 "Straight Waveguide" sch_x=107 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3947 N$7893 N$7894 "Straight Waveguide" sch_x=107 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3948 N$7895 N$7896 "Straight Waveguide" sch_x=107 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3949 N$7897 N$7898 "Straight Waveguide" sch_x=107 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3950 N$7899 N$7900 "Straight Waveguide" sch_x=107 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3951 N$7901 N$7902 "Straight Waveguide" sch_x=107 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3952 N$7903 N$7904 "Straight Waveguide" sch_x=107 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3953 N$7905 N$7906 "Straight Waveguide" sch_x=107 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3954 N$7907 N$7908 "Straight Waveguide" sch_x=107 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3955 N$7909 N$7910 "Straight Waveguide" sch_x=105 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3956 N$7911 N$7912 "Straight Waveguide" sch_x=105 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3957 N$7913 N$7914 "Straight Waveguide" sch_x=105 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3958 N$7915 N$7916 "Straight Waveguide" sch_x=105 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3959 N$7917 N$7918 "Straight Waveguide" sch_x=105 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3960 N$7919 N$7920 "Straight Waveguide" sch_x=105 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3961 N$7921 N$7922 "Straight Waveguide" sch_x=105 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3962 N$7923 N$7924 "Straight Waveguide" sch_x=105 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3963 N$7925 N$7926 "Straight Waveguide" sch_x=105 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3964 N$7927 N$7928 "Straight Waveguide" sch_x=105 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3965 N$7929 N$7930 "Straight Waveguide" sch_x=105 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3966 N$7931 N$7932 "Straight Waveguide" sch_x=105 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3967 N$7933 N$7934 "Straight Waveguide" sch_x=105 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3968 N$7935 N$7936 "Straight Waveguide" sch_x=105 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3969 N$7937 N$7938 "Straight Waveguide" sch_x=105 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3970 N$7939 N$7940 "Straight Waveguide" sch_x=105 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3971 N$7941 N$7942 "Straight Waveguide" sch_x=105 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3972 N$7943 N$7944 "Straight Waveguide" sch_x=105 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3973 N$7945 N$7946 "Straight Waveguide" sch_x=105 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3974 N$7947 N$7948 "Straight Waveguide" sch_x=105 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3975 N$7949 N$7950 "Straight Waveguide" sch_x=105 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3976 N$7951 N$7952 "Straight Waveguide" sch_x=105 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3977 N$7953 N$7954 "Straight Waveguide" sch_x=105 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3978 N$7955 N$7956 "Straight Waveguide" sch_x=105 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3979 N$7957 N$7958 "Straight Waveguide" sch_x=105 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3980 N$7959 N$7960 "Straight Waveguide" sch_x=105 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3981 N$7961 N$7962 "Straight Waveguide" sch_x=105 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3982 N$7963 N$7964 "Straight Waveguide" sch_x=105 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3983 N$7965 N$7966 "Straight Waveguide" sch_x=105 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3984 N$7967 N$7968 "Straight Waveguide" sch_x=105 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3985 N$7969 N$7970 "Straight Waveguide" sch_x=105 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3986 N$7971 N$7972 "Straight Waveguide" sch_x=105 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3987 N$7973 N$7974 "Straight Waveguide" sch_x=105 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3988 N$7975 N$7976 "Straight Waveguide" sch_x=105 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3989 N$7977 N$7978 "Straight Waveguide" sch_x=105 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3990 N$7979 N$7980 "Straight Waveguide" sch_x=105 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3991 N$7981 N$7982 "Straight Waveguide" sch_x=105 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3992 N$7983 N$7984 "Straight Waveguide" sch_x=105 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3993 N$7985 N$7986 "Straight Waveguide" sch_x=105 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3994 N$7987 N$7988 "Straight Waveguide" sch_x=105 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3995 N$7989 N$7990 "Straight Waveguide" sch_x=105 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3996 N$7991 N$7992 "Straight Waveguide" sch_x=105 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3997 N$7993 N$7994 "Straight Waveguide" sch_x=103 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3998 N$7995 N$7996 "Straight Waveguide" sch_x=103 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3999 N$7997 N$7998 "Straight Waveguide" sch_x=103 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4000 N$7999 N$8000 "Straight Waveguide" sch_x=103 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4001 N$8001 N$8002 "Straight Waveguide" sch_x=103 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4002 N$8003 N$8004 "Straight Waveguide" sch_x=103 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4003 N$8005 N$8006 "Straight Waveguide" sch_x=103 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4004 N$8007 N$8008 "Straight Waveguide" sch_x=103 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4005 N$8009 N$8010 "Straight Waveguide" sch_x=103 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4006 N$8011 N$8012 "Straight Waveguide" sch_x=103 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4007 N$8013 N$8014 "Straight Waveguide" sch_x=103 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4008 N$8015 N$8016 "Straight Waveguide" sch_x=103 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4009 N$8017 N$8018 "Straight Waveguide" sch_x=103 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4010 N$8019 N$8020 "Straight Waveguide" sch_x=103 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4011 N$8021 N$8022 "Straight Waveguide" sch_x=103 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4012 N$8023 N$8024 "Straight Waveguide" sch_x=103 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4013 N$8025 N$8026 "Straight Waveguide" sch_x=103 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4014 N$8027 N$8028 "Straight Waveguide" sch_x=103 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4015 N$8029 N$8030 "Straight Waveguide" sch_x=103 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4016 N$8031 N$8032 "Straight Waveguide" sch_x=103 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4017 N$8033 N$8034 "Straight Waveguide" sch_x=103 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4018 N$8035 N$8036 "Straight Waveguide" sch_x=103 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4019 N$8037 N$8038 "Straight Waveguide" sch_x=103 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4020 N$8039 N$8040 "Straight Waveguide" sch_x=103 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4021 N$8041 N$8042 "Straight Waveguide" sch_x=103 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4022 N$8043 N$8044 "Straight Waveguide" sch_x=103 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4023 N$8045 N$8046 "Straight Waveguide" sch_x=103 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4024 N$8047 N$8048 "Straight Waveguide" sch_x=103 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4025 N$8049 N$8050 "Straight Waveguide" sch_x=103 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4026 N$8051 N$8052 "Straight Waveguide" sch_x=103 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4027 N$8053 N$8054 "Straight Waveguide" sch_x=103 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4028 N$8055 N$8056 "Straight Waveguide" sch_x=103 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4029 N$8057 N$8058 "Straight Waveguide" sch_x=103 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4030 N$8059 N$8060 "Straight Waveguide" sch_x=103 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4031 N$8061 N$8062 "Straight Waveguide" sch_x=103 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4032 N$8063 N$8064 "Straight Waveguide" sch_x=103 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4033 N$8065 N$8066 "Straight Waveguide" sch_x=103 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4034 N$8067 N$8068 "Straight Waveguide" sch_x=103 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4035 N$8069 N$8070 "Straight Waveguide" sch_x=103 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4036 N$8071 N$8072 "Straight Waveguide" sch_x=103 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4037 N$8073 N$8074 "Straight Waveguide" sch_x=101 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4038 N$8075 N$8076 "Straight Waveguide" sch_x=101 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4039 N$8077 N$8078 "Straight Waveguide" sch_x=101 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4040 N$8079 N$8080 "Straight Waveguide" sch_x=101 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4041 N$8081 N$8082 "Straight Waveguide" sch_x=101 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4042 N$8083 N$8084 "Straight Waveguide" sch_x=101 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4043 N$8085 N$8086 "Straight Waveguide" sch_x=101 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4044 N$8087 N$8088 "Straight Waveguide" sch_x=101 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4045 N$8089 N$8090 "Straight Waveguide" sch_x=101 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4046 N$8091 N$8092 "Straight Waveguide" sch_x=101 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4047 N$8093 N$8094 "Straight Waveguide" sch_x=101 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4048 N$8095 N$8096 "Straight Waveguide" sch_x=101 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4049 N$8097 N$8098 "Straight Waveguide" sch_x=101 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4050 N$8099 N$8100 "Straight Waveguide" sch_x=101 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4051 N$8101 N$8102 "Straight Waveguide" sch_x=101 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4052 N$8103 N$8104 "Straight Waveguide" sch_x=101 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4053 N$8105 N$8106 "Straight Waveguide" sch_x=101 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4054 N$8107 N$8108 "Straight Waveguide" sch_x=101 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4055 N$8109 N$8110 "Straight Waveguide" sch_x=101 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4056 N$8111 N$8112 "Straight Waveguide" sch_x=101 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4057 N$8113 N$8114 "Straight Waveguide" sch_x=101 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4058 N$8115 N$8116 "Straight Waveguide" sch_x=101 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4059 N$8117 N$8118 "Straight Waveguide" sch_x=101 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4060 N$8119 N$8120 "Straight Waveguide" sch_x=101 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4061 N$8121 N$8122 "Straight Waveguide" sch_x=101 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4062 N$8123 N$8124 "Straight Waveguide" sch_x=101 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4063 N$8125 N$8126 "Straight Waveguide" sch_x=101 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4064 N$8127 N$8128 "Straight Waveguide" sch_x=101 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4065 N$8129 N$8130 "Straight Waveguide" sch_x=101 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4066 N$8131 N$8132 "Straight Waveguide" sch_x=101 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4067 N$8133 N$8134 "Straight Waveguide" sch_x=101 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4068 N$8135 N$8136 "Straight Waveguide" sch_x=101 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4069 N$8137 N$8138 "Straight Waveguide" sch_x=101 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4070 N$8139 N$8140 "Straight Waveguide" sch_x=101 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4071 N$8141 N$8142 "Straight Waveguide" sch_x=101 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4072 N$8143 N$8144 "Straight Waveguide" sch_x=101 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4073 N$8145 N$8146 "Straight Waveguide" sch_x=101 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4074 N$8147 N$8148 "Straight Waveguide" sch_x=101 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4075 N$8149 N$8150 "Straight Waveguide" sch_x=99 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4076 N$8151 N$8152 "Straight Waveguide" sch_x=99 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4077 N$8153 N$8154 "Straight Waveguide" sch_x=99 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4078 N$8155 N$8156 "Straight Waveguide" sch_x=99 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4079 N$8157 N$8158 "Straight Waveguide" sch_x=99 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4080 N$8159 N$8160 "Straight Waveguide" sch_x=99 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4081 N$8161 N$8162 "Straight Waveguide" sch_x=99 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4082 N$8163 N$8164 "Straight Waveguide" sch_x=99 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4083 N$8165 N$8166 "Straight Waveguide" sch_x=99 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4084 N$8167 N$8168 "Straight Waveguide" sch_x=99 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4085 N$8169 N$8170 "Straight Waveguide" sch_x=99 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4086 N$8171 N$8172 "Straight Waveguide" sch_x=99 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4087 N$8173 N$8174 "Straight Waveguide" sch_x=99 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4088 N$8175 N$8176 "Straight Waveguide" sch_x=99 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4089 N$8177 N$8178 "Straight Waveguide" sch_x=99 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4090 N$8179 N$8180 "Straight Waveguide" sch_x=99 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4091 N$8181 N$8182 "Straight Waveguide" sch_x=99 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4092 N$8183 N$8184 "Straight Waveguide" sch_x=99 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4093 N$8185 N$8186 "Straight Waveguide" sch_x=99 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4094 N$8187 N$8188 "Straight Waveguide" sch_x=99 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4095 N$8189 N$8190 "Straight Waveguide" sch_x=99 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4096 N$8191 N$8192 "Straight Waveguide" sch_x=99 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4097 N$8193 N$8194 "Straight Waveguide" sch_x=99 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4098 N$8195 N$8196 "Straight Waveguide" sch_x=99 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4099 N$8197 N$8198 "Straight Waveguide" sch_x=99 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4100 N$8199 N$8200 "Straight Waveguide" sch_x=99 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4101 N$8201 N$8202 "Straight Waveguide" sch_x=99 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4102 N$8203 N$8204 "Straight Waveguide" sch_x=99 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4103 N$8205 N$8206 "Straight Waveguide" sch_x=99 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4104 N$8207 N$8208 "Straight Waveguide" sch_x=99 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4105 N$8209 N$8210 "Straight Waveguide" sch_x=99 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4106 N$8211 N$8212 "Straight Waveguide" sch_x=99 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4107 N$8213 N$8214 "Straight Waveguide" sch_x=99 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4108 N$8215 N$8216 "Straight Waveguide" sch_x=99 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4109 N$8217 N$8218 "Straight Waveguide" sch_x=99 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4110 N$8219 N$8220 "Straight Waveguide" sch_x=99 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4111 N$8221 N$8222 "Straight Waveguide" sch_x=97 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4112 N$8223 N$8224 "Straight Waveguide" sch_x=97 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4113 N$8225 N$8226 "Straight Waveguide" sch_x=97 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4114 N$8227 N$8228 "Straight Waveguide" sch_x=97 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4115 N$8229 N$8230 "Straight Waveguide" sch_x=97 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4116 N$8231 N$8232 "Straight Waveguide" sch_x=97 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4117 N$8233 N$8234 "Straight Waveguide" sch_x=97 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4118 N$8235 N$8236 "Straight Waveguide" sch_x=97 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4119 N$8237 N$8238 "Straight Waveguide" sch_x=97 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4120 N$8239 N$8240 "Straight Waveguide" sch_x=97 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4121 N$8241 N$8242 "Straight Waveguide" sch_x=97 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4122 N$8243 N$8244 "Straight Waveguide" sch_x=97 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4123 N$8245 N$8246 "Straight Waveguide" sch_x=97 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4124 N$8247 N$8248 "Straight Waveguide" sch_x=97 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4125 N$8249 N$8250 "Straight Waveguide" sch_x=97 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4126 N$8251 N$8252 "Straight Waveguide" sch_x=97 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4127 N$8253 N$8254 "Straight Waveguide" sch_x=97 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4128 N$8255 N$8256 "Straight Waveguide" sch_x=97 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4129 N$8257 N$8258 "Straight Waveguide" sch_x=97 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4130 N$8259 N$8260 "Straight Waveguide" sch_x=97 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4131 N$8261 N$8262 "Straight Waveguide" sch_x=97 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4132 N$8263 N$8264 "Straight Waveguide" sch_x=97 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4133 N$8265 N$8266 "Straight Waveguide" sch_x=97 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4134 N$8267 N$8268 "Straight Waveguide" sch_x=97 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4135 N$8269 N$8270 "Straight Waveguide" sch_x=97 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4136 N$8271 N$8272 "Straight Waveguide" sch_x=97 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4137 N$8273 N$8274 "Straight Waveguide" sch_x=97 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4138 N$8275 N$8276 "Straight Waveguide" sch_x=97 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4139 N$8277 N$8278 "Straight Waveguide" sch_x=97 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4140 N$8279 N$8280 "Straight Waveguide" sch_x=97 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4141 N$8281 N$8282 "Straight Waveguide" sch_x=97 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4142 N$8283 N$8284 "Straight Waveguide" sch_x=97 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4143 N$8285 N$8286 "Straight Waveguide" sch_x=97 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4144 N$8287 N$8288 "Straight Waveguide" sch_x=97 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4145 N$8289 N$8290 "Straight Waveguide" sch_x=95 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4146 N$8291 N$8292 "Straight Waveguide" sch_x=95 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4147 N$8293 N$8294 "Straight Waveguide" sch_x=95 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4148 N$8295 N$8296 "Straight Waveguide" sch_x=95 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4149 N$8297 N$8298 "Straight Waveguide" sch_x=95 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4150 N$8299 N$8300 "Straight Waveguide" sch_x=95 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4151 N$8301 N$8302 "Straight Waveguide" sch_x=95 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4152 N$8303 N$8304 "Straight Waveguide" sch_x=95 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4153 N$8305 N$8306 "Straight Waveguide" sch_x=95 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4154 N$8307 N$8308 "Straight Waveguide" sch_x=95 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4155 N$8309 N$8310 "Straight Waveguide" sch_x=95 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4156 N$8311 N$8312 "Straight Waveguide" sch_x=95 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4157 N$8313 N$8314 "Straight Waveguide" sch_x=95 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4158 N$8315 N$8316 "Straight Waveguide" sch_x=95 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4159 N$8317 N$8318 "Straight Waveguide" sch_x=95 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4160 N$8319 N$8320 "Straight Waveguide" sch_x=95 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4161 N$8321 N$8322 "Straight Waveguide" sch_x=95 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4162 N$8323 N$8324 "Straight Waveguide" sch_x=95 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4163 N$8325 N$8326 "Straight Waveguide" sch_x=95 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4164 N$8327 N$8328 "Straight Waveguide" sch_x=95 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4165 N$8329 N$8330 "Straight Waveguide" sch_x=95 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4166 N$8331 N$8332 "Straight Waveguide" sch_x=95 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4167 N$8333 N$8334 "Straight Waveguide" sch_x=95 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4168 N$8335 N$8336 "Straight Waveguide" sch_x=95 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4169 N$8337 N$8338 "Straight Waveguide" sch_x=95 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4170 N$8339 N$8340 "Straight Waveguide" sch_x=95 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4171 N$8341 N$8342 "Straight Waveguide" sch_x=95 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4172 N$8343 N$8344 "Straight Waveguide" sch_x=95 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4173 N$8345 N$8346 "Straight Waveguide" sch_x=95 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4174 N$8347 N$8348 "Straight Waveguide" sch_x=95 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4175 N$8349 N$8350 "Straight Waveguide" sch_x=95 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4176 N$8351 N$8352 "Straight Waveguide" sch_x=95 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4177 N$8353 N$8354 "Straight Waveguide" sch_x=93 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4178 N$8355 N$8356 "Straight Waveguide" sch_x=93 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4179 N$8357 N$8358 "Straight Waveguide" sch_x=93 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4180 N$8359 N$8360 "Straight Waveguide" sch_x=93 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4181 N$8361 N$8362 "Straight Waveguide" sch_x=93 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4182 N$8363 N$8364 "Straight Waveguide" sch_x=93 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4183 N$8365 N$8366 "Straight Waveguide" sch_x=93 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4184 N$8367 N$8368 "Straight Waveguide" sch_x=93 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4185 N$8369 N$8370 "Straight Waveguide" sch_x=93 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4186 N$8371 N$8372 "Straight Waveguide" sch_x=93 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4187 N$8373 N$8374 "Straight Waveguide" sch_x=93 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4188 N$8375 N$8376 "Straight Waveguide" sch_x=93 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4189 N$8377 N$8378 "Straight Waveguide" sch_x=93 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4190 N$8379 N$8380 "Straight Waveguide" sch_x=93 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4191 N$8381 N$8382 "Straight Waveguide" sch_x=93 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4192 N$8383 N$8384 "Straight Waveguide" sch_x=93 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4193 N$8385 N$8386 "Straight Waveguide" sch_x=93 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4194 N$8387 N$8388 "Straight Waveguide" sch_x=93 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4195 N$8389 N$8390 "Straight Waveguide" sch_x=93 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4196 N$8391 N$8392 "Straight Waveguide" sch_x=93 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4197 N$8393 N$8394 "Straight Waveguide" sch_x=93 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4198 N$8395 N$8396 "Straight Waveguide" sch_x=93 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4199 N$8397 N$8398 "Straight Waveguide" sch_x=93 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4200 N$8399 N$8400 "Straight Waveguide" sch_x=93 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4201 N$8401 N$8402 "Straight Waveguide" sch_x=93 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4202 N$8403 N$8404 "Straight Waveguide" sch_x=93 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4203 N$8405 N$8406 "Straight Waveguide" sch_x=93 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4204 N$8407 N$8408 "Straight Waveguide" sch_x=93 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4205 N$8409 N$8410 "Straight Waveguide" sch_x=93 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4206 N$8411 N$8412 "Straight Waveguide" sch_x=93 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4207 N$8413 N$8414 "Straight Waveguide" sch_x=91 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4208 N$8415 N$8416 "Straight Waveguide" sch_x=91 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4209 N$8417 N$8418 "Straight Waveguide" sch_x=91 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4210 N$8419 N$8420 "Straight Waveguide" sch_x=91 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4211 N$8421 N$8422 "Straight Waveguide" sch_x=91 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4212 N$8423 N$8424 "Straight Waveguide" sch_x=91 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4213 N$8425 N$8426 "Straight Waveguide" sch_x=91 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4214 N$8427 N$8428 "Straight Waveguide" sch_x=91 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4215 N$8429 N$8430 "Straight Waveguide" sch_x=91 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4216 N$8431 N$8432 "Straight Waveguide" sch_x=91 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4217 N$8433 N$8434 "Straight Waveguide" sch_x=91 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4218 N$8435 N$8436 "Straight Waveguide" sch_x=91 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4219 N$8437 N$8438 "Straight Waveguide" sch_x=91 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4220 N$8439 N$8440 "Straight Waveguide" sch_x=91 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4221 N$8441 N$8442 "Straight Waveguide" sch_x=91 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4222 N$8443 N$8444 "Straight Waveguide" sch_x=91 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4223 N$8445 N$8446 "Straight Waveguide" sch_x=91 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4224 N$8447 N$8448 "Straight Waveguide" sch_x=91 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4225 N$8449 N$8450 "Straight Waveguide" sch_x=91 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4226 N$8451 N$8452 "Straight Waveguide" sch_x=91 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4227 N$8453 N$8454 "Straight Waveguide" sch_x=91 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4228 N$8455 N$8456 "Straight Waveguide" sch_x=91 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4229 N$8457 N$8458 "Straight Waveguide" sch_x=91 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4230 N$8459 N$8460 "Straight Waveguide" sch_x=91 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4231 N$8461 N$8462 "Straight Waveguide" sch_x=91 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4232 N$8463 N$8464 "Straight Waveguide" sch_x=91 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4233 N$8465 N$8466 "Straight Waveguide" sch_x=91 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4234 N$8467 N$8468 "Straight Waveguide" sch_x=91 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4235 N$8469 N$8470 "Straight Waveguide" sch_x=89 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4236 N$8471 N$8472 "Straight Waveguide" sch_x=89 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4237 N$8473 N$8474 "Straight Waveguide" sch_x=89 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4238 N$8475 N$8476 "Straight Waveguide" sch_x=89 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4239 N$8477 N$8478 "Straight Waveguide" sch_x=89 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4240 N$8479 N$8480 "Straight Waveguide" sch_x=89 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4241 N$8481 N$8482 "Straight Waveguide" sch_x=89 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4242 N$8483 N$8484 "Straight Waveguide" sch_x=89 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4243 N$8485 N$8486 "Straight Waveguide" sch_x=89 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4244 N$8487 N$8488 "Straight Waveguide" sch_x=89 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4245 N$8489 N$8490 "Straight Waveguide" sch_x=89 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4246 N$8491 N$8492 "Straight Waveguide" sch_x=89 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4247 N$8493 N$8494 "Straight Waveguide" sch_x=89 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4248 N$8495 N$8496 "Straight Waveguide" sch_x=89 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4249 N$8497 N$8498 "Straight Waveguide" sch_x=89 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4250 N$8499 N$8500 "Straight Waveguide" sch_x=89 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4251 N$8501 N$8502 "Straight Waveguide" sch_x=89 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4252 N$8503 N$8504 "Straight Waveguide" sch_x=89 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4253 N$8505 N$8506 "Straight Waveguide" sch_x=89 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4254 N$8507 N$8508 "Straight Waveguide" sch_x=89 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4255 N$8509 N$8510 "Straight Waveguide" sch_x=89 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4256 N$8511 N$8512 "Straight Waveguide" sch_x=89 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4257 N$8513 N$8514 "Straight Waveguide" sch_x=89 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4258 N$8515 N$8516 "Straight Waveguide" sch_x=89 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4259 N$8517 N$8518 "Straight Waveguide" sch_x=89 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4260 N$8519 N$8520 "Straight Waveguide" sch_x=89 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4261 N$8521 N$8522 "Straight Waveguide" sch_x=87 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4262 N$8523 N$8524 "Straight Waveguide" sch_x=87 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4263 N$8525 N$8526 "Straight Waveguide" sch_x=87 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4264 N$8527 N$8528 "Straight Waveguide" sch_x=87 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4265 N$8529 N$8530 "Straight Waveguide" sch_x=87 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4266 N$8531 N$8532 "Straight Waveguide" sch_x=87 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4267 N$8533 N$8534 "Straight Waveguide" sch_x=87 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4268 N$8535 N$8536 "Straight Waveguide" sch_x=87 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4269 N$8537 N$8538 "Straight Waveguide" sch_x=87 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4270 N$8539 N$8540 "Straight Waveguide" sch_x=87 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4271 N$8541 N$8542 "Straight Waveguide" sch_x=87 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4272 N$8543 N$8544 "Straight Waveguide" sch_x=87 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4273 N$8545 N$8546 "Straight Waveguide" sch_x=87 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4274 N$8547 N$8548 "Straight Waveguide" sch_x=87 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4275 N$8549 N$8550 "Straight Waveguide" sch_x=87 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4276 N$8551 N$8552 "Straight Waveguide" sch_x=87 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4277 N$8553 N$8554 "Straight Waveguide" sch_x=87 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4278 N$8555 N$8556 "Straight Waveguide" sch_x=87 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4279 N$8557 N$8558 "Straight Waveguide" sch_x=87 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4280 N$8559 N$8560 "Straight Waveguide" sch_x=87 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4281 N$8561 N$8562 "Straight Waveguide" sch_x=87 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4282 N$8563 N$8564 "Straight Waveguide" sch_x=87 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4283 N$8565 N$8566 "Straight Waveguide" sch_x=87 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4284 N$8567 N$8568 "Straight Waveguide" sch_x=87 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4285 N$8569 N$8570 "Straight Waveguide" sch_x=85 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4286 N$8571 N$8572 "Straight Waveguide" sch_x=85 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4287 N$8573 N$8574 "Straight Waveguide" sch_x=85 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4288 N$8575 N$8576 "Straight Waveguide" sch_x=85 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4289 N$8577 N$8578 "Straight Waveguide" sch_x=85 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4290 N$8579 N$8580 "Straight Waveguide" sch_x=85 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4291 N$8581 N$8582 "Straight Waveguide" sch_x=85 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4292 N$8583 N$8584 "Straight Waveguide" sch_x=85 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4293 N$8585 N$8586 "Straight Waveguide" sch_x=85 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4294 N$8587 N$8588 "Straight Waveguide" sch_x=85 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4295 N$8589 N$8590 "Straight Waveguide" sch_x=85 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4296 N$8591 N$8592 "Straight Waveguide" sch_x=85 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4297 N$8593 N$8594 "Straight Waveguide" sch_x=85 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4298 N$8595 N$8596 "Straight Waveguide" sch_x=85 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4299 N$8597 N$8598 "Straight Waveguide" sch_x=85 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4300 N$8599 N$8600 "Straight Waveguide" sch_x=85 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4301 N$8601 N$8602 "Straight Waveguide" sch_x=85 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4302 N$8603 N$8604 "Straight Waveguide" sch_x=85 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4303 N$8605 N$8606 "Straight Waveguide" sch_x=85 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4304 N$8607 N$8608 "Straight Waveguide" sch_x=85 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4305 N$8609 N$8610 "Straight Waveguide" sch_x=85 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4306 N$8611 N$8612 "Straight Waveguide" sch_x=85 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4307 N$8613 N$8614 "Straight Waveguide" sch_x=83 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4308 N$8615 N$8616 "Straight Waveguide" sch_x=83 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4309 N$8617 N$8618 "Straight Waveguide" sch_x=83 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4310 N$8619 N$8620 "Straight Waveguide" sch_x=83 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4311 N$8621 N$8622 "Straight Waveguide" sch_x=83 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4312 N$8623 N$8624 "Straight Waveguide" sch_x=83 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4313 N$8625 N$8626 "Straight Waveguide" sch_x=83 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4314 N$8627 N$8628 "Straight Waveguide" sch_x=83 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4315 N$8629 N$8630 "Straight Waveguide" sch_x=83 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4316 N$8631 N$8632 "Straight Waveguide" sch_x=83 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4317 N$8633 N$8634 "Straight Waveguide" sch_x=83 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4318 N$8635 N$8636 "Straight Waveguide" sch_x=83 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4319 N$8637 N$8638 "Straight Waveguide" sch_x=83 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4320 N$8639 N$8640 "Straight Waveguide" sch_x=83 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4321 N$8641 N$8642 "Straight Waveguide" sch_x=83 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4322 N$8643 N$8644 "Straight Waveguide" sch_x=83 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4323 N$8645 N$8646 "Straight Waveguide" sch_x=83 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4324 N$8647 N$8648 "Straight Waveguide" sch_x=83 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4325 N$8649 N$8650 "Straight Waveguide" sch_x=83 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4326 N$8651 N$8652 "Straight Waveguide" sch_x=83 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4327 N$8653 N$8654 "Straight Waveguide" sch_x=81 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4328 N$8655 N$8656 "Straight Waveguide" sch_x=81 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4329 N$8657 N$8658 "Straight Waveguide" sch_x=81 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4330 N$8659 N$8660 "Straight Waveguide" sch_x=81 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4331 N$8661 N$8662 "Straight Waveguide" sch_x=81 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4332 N$8663 N$8664 "Straight Waveguide" sch_x=81 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4333 N$8665 N$8666 "Straight Waveguide" sch_x=81 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4334 N$8667 N$8668 "Straight Waveguide" sch_x=81 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4335 N$8669 N$8670 "Straight Waveguide" sch_x=81 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4336 N$8671 N$8672 "Straight Waveguide" sch_x=81 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4337 N$8673 N$8674 "Straight Waveguide" sch_x=81 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4338 N$8675 N$8676 "Straight Waveguide" sch_x=81 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4339 N$8677 N$8678 "Straight Waveguide" sch_x=81 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4340 N$8679 N$8680 "Straight Waveguide" sch_x=81 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4341 N$8681 N$8682 "Straight Waveguide" sch_x=81 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4342 N$8683 N$8684 "Straight Waveguide" sch_x=81 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4343 N$8685 N$8686 "Straight Waveguide" sch_x=81 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4344 N$8687 N$8688 "Straight Waveguide" sch_x=81 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4345 N$8689 N$8690 "Straight Waveguide" sch_x=79 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4346 N$8691 N$8692 "Straight Waveguide" sch_x=79 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4347 N$8693 N$8694 "Straight Waveguide" sch_x=79 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4348 N$8695 N$8696 "Straight Waveguide" sch_x=79 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4349 N$8697 N$8698 "Straight Waveguide" sch_x=79 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4350 N$8699 N$8700 "Straight Waveguide" sch_x=79 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4351 N$8701 N$8702 "Straight Waveguide" sch_x=79 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4352 N$8703 N$8704 "Straight Waveguide" sch_x=79 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4353 N$8705 N$8706 "Straight Waveguide" sch_x=79 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4354 N$8707 N$8708 "Straight Waveguide" sch_x=79 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4355 N$8709 N$8710 "Straight Waveguide" sch_x=79 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4356 N$8711 N$8712 "Straight Waveguide" sch_x=79 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4357 N$8713 N$8714 "Straight Waveguide" sch_x=79 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4358 N$8715 N$8716 "Straight Waveguide" sch_x=79 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4359 N$8717 N$8718 "Straight Waveguide" sch_x=79 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4360 N$8719 N$8720 "Straight Waveguide" sch_x=79 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4361 N$8721 N$8722 "Straight Waveguide" sch_x=77 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4362 N$8723 N$8724 "Straight Waveguide" sch_x=77 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4363 N$8725 N$8726 "Straight Waveguide" sch_x=77 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4364 N$8727 N$8728 "Straight Waveguide" sch_x=77 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4365 N$8729 N$8730 "Straight Waveguide" sch_x=77 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4366 N$8731 N$8732 "Straight Waveguide" sch_x=77 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4367 N$8733 N$8734 "Straight Waveguide" sch_x=77 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4368 N$8735 N$8736 "Straight Waveguide" sch_x=77 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4369 N$8737 N$8738 "Straight Waveguide" sch_x=77 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4370 N$8739 N$8740 "Straight Waveguide" sch_x=77 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4371 N$8741 N$8742 "Straight Waveguide" sch_x=77 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4372 N$8743 N$8744 "Straight Waveguide" sch_x=77 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4373 N$8745 N$8746 "Straight Waveguide" sch_x=77 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4374 N$8747 N$8748 "Straight Waveguide" sch_x=77 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4375 N$8749 N$8750 "Straight Waveguide" sch_x=75 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4376 N$8751 N$8752 "Straight Waveguide" sch_x=75 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4377 N$8753 N$8754 "Straight Waveguide" sch_x=75 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4378 N$8755 N$8756 "Straight Waveguide" sch_x=75 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4379 N$8757 N$8758 "Straight Waveguide" sch_x=75 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4380 N$8759 N$8760 "Straight Waveguide" sch_x=75 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4381 N$8761 N$8762 "Straight Waveguide" sch_x=75 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4382 N$8763 N$8764 "Straight Waveguide" sch_x=75 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4383 N$8765 N$8766 "Straight Waveguide" sch_x=75 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4384 N$8767 N$8768 "Straight Waveguide" sch_x=75 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4385 N$8769 N$8770 "Straight Waveguide" sch_x=75 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4386 N$8771 N$8772 "Straight Waveguide" sch_x=75 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4387 N$8773 N$8774 "Straight Waveguide" sch_x=73 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4388 N$8775 N$8776 "Straight Waveguide" sch_x=73 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4389 N$8777 N$8778 "Straight Waveguide" sch_x=73 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4390 N$8779 N$8780 "Straight Waveguide" sch_x=73 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4391 N$8781 N$8782 "Straight Waveguide" sch_x=73 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4392 N$8783 N$8784 "Straight Waveguide" sch_x=73 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4393 N$8785 N$8786 "Straight Waveguide" sch_x=73 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4394 N$8787 N$8788 "Straight Waveguide" sch_x=73 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4395 N$8789 N$8790 "Straight Waveguide" sch_x=73 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4396 N$8791 N$8792 "Straight Waveguide" sch_x=73 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4397 N$8793 N$8794 "Straight Waveguide" sch_x=71 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4398 N$8795 N$8796 "Straight Waveguide" sch_x=71 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4399 N$8797 N$8798 "Straight Waveguide" sch_x=71 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4400 N$8799 N$8800 "Straight Waveguide" sch_x=71 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4401 N$8801 N$8802 "Straight Waveguide" sch_x=71 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4402 N$8803 N$8804 "Straight Waveguide" sch_x=71 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4403 N$8805 N$8806 "Straight Waveguide" sch_x=71 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4404 N$8807 N$8808 "Straight Waveguide" sch_x=71 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4405 N$8809 N$8810 "Straight Waveguide" sch_x=69 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4406 N$8811 N$8812 "Straight Waveguide" sch_x=69 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4407 N$8813 N$8814 "Straight Waveguide" sch_x=69 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4408 N$8815 N$8816 "Straight Waveguide" sch_x=69 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4409 N$8817 N$8818 "Straight Waveguide" sch_x=69 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4410 N$8819 N$8820 "Straight Waveguide" sch_x=69 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4411 N$8821 N$8822 "Straight Waveguide" sch_x=67 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4412 N$8823 N$8824 "Straight Waveguide" sch_x=67 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4413 N$8825 N$8826 "Straight Waveguide" sch_x=67 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4414 N$8827 N$8828 "Straight Waveguide" sch_x=67 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4415 N$8829 N$8830 "Straight Waveguide" sch_x=65 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4416 N$8831 N$8832 "Straight Waveguide" sch_x=65 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4417 N$8834 N$8833 "Straight Waveguide" sch_x=93 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4418 N$8836 N$8835 "Straight Waveguide" sch_x=92 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4419 N$8838 N$8837 "Straight Waveguide" sch_x=91 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4420 N$8840 N$8839 "Straight Waveguide" sch_x=90 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4421 N$8842 N$8841 "Straight Waveguide" sch_x=89 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4422 N$8844 N$8843 "Straight Waveguide" sch_x=88 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4423 N$8846 N$8845 "Straight Waveguide" sch_x=87 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4424 N$8848 N$8847 "Straight Waveguide" sch_x=86 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4425 N$8850 N$8849 "Straight Waveguide" sch_x=85 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4426 N$8852 N$8851 "Straight Waveguide" sch_x=84 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4427 N$8854 N$8853 "Straight Waveguide" sch_x=83 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4428 N$8856 N$8855 "Straight Waveguide" sch_x=82 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4429 N$8858 N$8857 "Straight Waveguide" sch_x=81 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4430 N$8860 N$8859 "Straight Waveguide" sch_x=80 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4431 N$8862 N$8861 "Straight Waveguide" sch_x=79 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4432 N$8864 N$8863 "Straight Waveguide" sch_x=78 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4433 N$8866 N$8865 "Straight Waveguide" sch_x=77 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4434 N$8868 N$8867 "Straight Waveguide" sch_x=76 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4435 N$8870 N$8869 "Straight Waveguide" sch_x=75 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4436 N$8872 N$8871 "Straight Waveguide" sch_x=74 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4437 N$8874 N$8873 "Straight Waveguide" sch_x=73 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4438 N$8876 N$8875 "Straight Waveguide" sch_x=72 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4439 N$8878 N$8877 "Straight Waveguide" sch_x=71 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4440 N$8880 N$8879 "Straight Waveguide" sch_x=70 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4441 N$8882 N$8881 "Straight Waveguide" sch_x=69 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4442 N$8884 N$8883 "Straight Waveguide" sch_x=68 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4443 N$8886 N$8885 "Straight Waveguide" sch_x=67 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4444 N$8888 N$8887 "Straight Waveguide" sch_x=66 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4445 N$8890 N$8889 "Straight Waveguide" sch_x=65 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4446 N$8892 N$8891 "Straight Waveguide" sch_x=64 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4447 N$8894 N$8893 "Straight Waveguide" sch_x=63 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4448 N$8896 N$8895 "Straight Waveguide" sch_x=63 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4449 N$8898 N$8897 "Straight Waveguide" sch_x=64 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4450 N$8900 N$8899 "Straight Waveguide" sch_x=65 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4451 N$8902 N$8901 "Straight Waveguide" sch_x=66 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4452 N$8904 N$8903 "Straight Waveguide" sch_x=67 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4453 N$8906 N$8905 "Straight Waveguide" sch_x=68 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4454 N$8908 N$8907 "Straight Waveguide" sch_x=69 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4455 N$8910 N$8909 "Straight Waveguide" sch_x=70 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4456 N$8912 N$8911 "Straight Waveguide" sch_x=71 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4457 N$8914 N$8913 "Straight Waveguide" sch_x=72 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4458 N$8916 N$8915 "Straight Waveguide" sch_x=73 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4459 N$8918 N$8917 "Straight Waveguide" sch_x=74 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4460 N$8920 N$8919 "Straight Waveguide" sch_x=75 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4461 N$8922 N$8921 "Straight Waveguide" sch_x=76 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4462 N$8924 N$8923 "Straight Waveguide" sch_x=77 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4463 N$8926 N$8925 "Straight Waveguide" sch_x=78 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4464 N$8928 N$8927 "Straight Waveguide" sch_x=79 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4465 N$8930 N$8929 "Straight Waveguide" sch_x=80 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4466 N$8932 N$8931 "Straight Waveguide" sch_x=81 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4467 N$8934 N$8933 "Straight Waveguide" sch_x=82 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4468 N$8936 N$8935 "Straight Waveguide" sch_x=83 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4469 N$8938 N$8937 "Straight Waveguide" sch_x=84 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4470 N$8940 N$8939 "Straight Waveguide" sch_x=85 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4471 N$8942 N$8941 "Straight Waveguide" sch_x=86 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4472 N$8944 N$8943 "Straight Waveguide" sch_x=87 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4473 N$8946 N$8945 "Straight Waveguide" sch_x=88 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4474 N$8948 N$8947 "Straight Waveguide" sch_x=89 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4475 N$8950 N$8949 "Straight Waveguide" sch_x=90 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4476 N$8952 N$8951 "Straight Waveguide" sch_x=91 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4477 N$8954 N$8953 "Straight Waveguide" sch_x=92 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4478 N$8956 N$8955 "Straight Waveguide" sch_x=93 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4479 N$8958 N$8957 "Straight Waveguide" sch_x=94 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4480 N$8960 N$8959 "Straight Waveguide" sch_x=94 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4481 N$8961 N$8962 "Straight Waveguide" sch_x=-4 sch_y=-0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4482 N$8963 N$8964 "Straight Waveguide" sch_x=-5 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4483 N$8965 N$8966 "Straight Waveguide" sch_x=-5 sch_y=-2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4484 N$8967 N$8968 "Straight Waveguide" sch_x=-3 sch_y=-1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4485 N$8969 N$8970 "Straight Waveguide" sch_x=-3 sch_y=-2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4486 N$8971 N$8972 "Straight Waveguide" sch_x=-4 sch_y=-3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4487 N$8973 N$8974 "Straight Waveguide" sch_x=0 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4488 N$8975 N$8976 "Straight Waveguide" sch_x=-1 sch_y=-0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4489 N$8977 N$8978 "Straight Waveguide" sch_x=-1 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4490 N$8979 N$8980 "Straight Waveguide" sch_x=1 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4491 N$8981 N$8982 "Straight Waveguide" sch_x=1 sch_y=-0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4492 N$8983 N$8984 "Straight Waveguide" sch_x=0 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4493 N$8985 N$8986 "Straight Waveguide" sch_x=0 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4494 N$8987 N$8988 "Straight Waveguide" sch_x=-1 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4495 N$8989 N$8990 "Straight Waveguide" sch_x=-1 sch_y=-3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4496 N$8991 N$8992 "Straight Waveguide" sch_x=1 sch_y=-3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4497 N$8993 N$8994 "Straight Waveguide" sch_x=1 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4498 N$8995 N$8996 "Straight Waveguide" sch_x=0 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4499 N$8997 N$8998 "Straight Waveguide" sch_x=4 sch_y=-0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4500 N$8999 N$9000 "Straight Waveguide" sch_x=3 sch_y=-1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4501 N$9001 N$9002 "Straight Waveguide" sch_x=3 sch_y=-2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4502 N$9003 N$9004 "Straight Waveguide" sch_x=5 sch_y=-2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4503 N$9005 N$9006 "Straight Waveguide" sch_x=5 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4504 N$9007 N$9008 "Straight Waveguide" sch_x=4 sch_y=-3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4505 N$9009 N$9010 "Straight Waveguide" sch_x=-4 sch_y=-4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4506 N$9011 N$9012 "Straight Waveguide" sch_x=-5 sch_y=-5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4507 N$9013 N$9014 "Straight Waveguide" sch_x=-5 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4508 N$9015 N$9016 "Straight Waveguide" sch_x=-3 sch_y=-5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4509 N$9017 N$9018 "Straight Waveguide" sch_x=-3 sch_y=-6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4510 N$9019 N$9020 "Straight Waveguide" sch_x=-4 sch_y=-7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4511 N$9021 N$9022 "Straight Waveguide" sch_x=0 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4512 N$9023 N$9024 "Straight Waveguide" sch_x=-1 sch_y=-4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4513 N$9025 N$9026 "Straight Waveguide" sch_x=-1 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4514 N$9027 N$9028 "Straight Waveguide" sch_x=1 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4515 N$9029 N$9030 "Straight Waveguide" sch_x=1 sch_y=-4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4516 N$9031 N$9032 "Straight Waveguide" sch_x=0 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4517 N$9033 N$9034 "Straight Waveguide" sch_x=0 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4518 N$9035 N$9036 "Straight Waveguide" sch_x=-1 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4519 N$9037 N$9038 "Straight Waveguide" sch_x=-1 sch_y=-7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4520 N$9039 N$9040 "Straight Waveguide" sch_x=1 sch_y=-7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4521 N$9041 N$9042 "Straight Waveguide" sch_x=1 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4522 N$9043 N$9044 "Straight Waveguide" sch_x=0 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4523 N$9045 N$9046 "Straight Waveguide" sch_x=4 sch_y=-4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4524 N$9047 N$9048 "Straight Waveguide" sch_x=3 sch_y=-5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4525 N$9049 N$9050 "Straight Waveguide" sch_x=3 sch_y=-6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4526 N$9051 N$9052 "Straight Waveguide" sch_x=5 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4527 N$9053 N$9054 "Straight Waveguide" sch_x=5 sch_y=-5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4528 N$9055 N$9056 "Straight Waveguide" sch_x=4 sch_y=-7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4529 N$9058 N$9057 "Straight Waveguide" sch_x=-13 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4530 N$9060 N$9059 "Straight Waveguide" sch_x=-13 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4531 N$9062 N$9061 "Straight Waveguide" sch_x=-13 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4532 N$9064 N$9063 "Straight Waveguide" sch_x=-13 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4533 N$9066 N$9065 "Straight Waveguide" sch_x=-13 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4534 N$9068 N$9067 "Straight Waveguide" sch_x=-13 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4535 N$9070 N$9069 "Straight Waveguide" sch_x=-11 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4536 N$9072 N$9071 "Straight Waveguide" sch_x=-11 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4537 N$9074 N$9073 "Straight Waveguide" sch_x=-11 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4538 N$9076 N$9075 "Straight Waveguide" sch_x=-11 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4539 N$9078 N$9077 "Straight Waveguide" sch_x=-9 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4540 N$9080 N$9079 "Straight Waveguide" sch_x=-9 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4541 N$9081 N$9082 "Straight Waveguide" sch_x=-9 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4542 N$9083 N$9084 "Straight Waveguide" sch_x=-8 sch_y=-2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4543 N$9085 N$9086 "Straight Waveguide" sch_x=-7 sch_y=-3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4544 N$9087 N$9088 "Straight Waveguide" sch_x=-7 sch_y=-4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4545 N$9089 N$9090 "Straight Waveguide" sch_x=-8 sch_y=-5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4546 N$9091 N$9092 "Straight Waveguide" sch_x=-9 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4547 N$9093 N$9094 "Straight Waveguide" sch_x=-10 sch_y=-1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4548 N$9095 N$9096 "Straight Waveguide" sch_x=-10 sch_y=-6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4549 N$9097 N$9098 "Straight Waveguide" sch_x=13 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4550 N$9099 N$9100 "Straight Waveguide" sch_x=13 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4551 N$9101 N$9102 "Straight Waveguide" sch_x=13 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4552 N$9103 N$9104 "Straight Waveguide" sch_x=13 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4553 N$9105 N$9106 "Straight Waveguide" sch_x=13 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4554 N$9107 N$9108 "Straight Waveguide" sch_x=13 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4555 N$9109 N$9110 "Straight Waveguide" sch_x=11 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4556 N$9111 N$9112 "Straight Waveguide" sch_x=11 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4557 N$9113 N$9114 "Straight Waveguide" sch_x=11 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4558 N$9115 N$9116 "Straight Waveguide" sch_x=11 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4559 N$9117 N$9118 "Straight Waveguide" sch_x=9 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4560 N$9119 N$9120 "Straight Waveguide" sch_x=9 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4561 N$9122 N$9121 "Straight Waveguide" sch_x=9 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4562 N$9124 N$9123 "Straight Waveguide" sch_x=8 sch_y=-2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4563 N$9126 N$9125 "Straight Waveguide" sch_x=7 sch_y=-3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4564 N$9128 N$9127 "Straight Waveguide" sch_x=7 sch_y=-4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4565 N$9130 N$9129 "Straight Waveguide" sch_x=8 sch_y=-5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4566 N$9132 N$9131 "Straight Waveguide" sch_x=9 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4567 N$9134 N$9133 "Straight Waveguide" sch_x=10 sch_y=-1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4568 N$9136 N$9135 "Straight Waveguide" sch_x=10 sch_y=-6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4569 N$9137 N$9138 "Straight Waveguide" sch_x=-4 sch_y=-8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4570 N$9139 N$9140 "Straight Waveguide" sch_x=-5 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4571 N$9141 N$9142 "Straight Waveguide" sch_x=-5 sch_y=-10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4572 N$9143 N$9144 "Straight Waveguide" sch_x=-3 sch_y=-9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4573 N$9145 N$9146 "Straight Waveguide" sch_x=-3 sch_y=-10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4574 N$9147 N$9148 "Straight Waveguide" sch_x=-4 sch_y=-11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4575 N$9149 N$9150 "Straight Waveguide" sch_x=0 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4576 N$9151 N$9152 "Straight Waveguide" sch_x=-1 sch_y=-8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4577 N$9153 N$9154 "Straight Waveguide" sch_x=-1 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4578 N$9155 N$9156 "Straight Waveguide" sch_x=1 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4579 N$9157 N$9158 "Straight Waveguide" sch_x=1 sch_y=-8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4580 N$9159 N$9160 "Straight Waveguide" sch_x=0 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4581 N$9161 N$9162 "Straight Waveguide" sch_x=0 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4582 N$9163 N$9164 "Straight Waveguide" sch_x=-1 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4583 N$9165 N$9166 "Straight Waveguide" sch_x=-1 sch_y=-11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4584 N$9167 N$9168 "Straight Waveguide" sch_x=1 sch_y=-11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4585 N$9169 N$9170 "Straight Waveguide" sch_x=1 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4586 N$9171 N$9172 "Straight Waveguide" sch_x=0 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4587 N$9173 N$9174 "Straight Waveguide" sch_x=4 sch_y=-8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4588 N$9175 N$9176 "Straight Waveguide" sch_x=3 sch_y=-9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4589 N$9177 N$9178 "Straight Waveguide" sch_x=3 sch_y=-10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4590 N$9179 N$9180 "Straight Waveguide" sch_x=5 sch_y=-10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4591 N$9181 N$9182 "Straight Waveguide" sch_x=5 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4592 N$9183 N$9184 "Straight Waveguide" sch_x=4 sch_y=-11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4593 N$9185 N$9186 "Straight Waveguide" sch_x=-4 sch_y=-12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4594 N$9187 N$9188 "Straight Waveguide" sch_x=-5 sch_y=-13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4595 N$9189 N$9190 "Straight Waveguide" sch_x=-5 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4596 N$9191 N$9192 "Straight Waveguide" sch_x=-3 sch_y=-13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4597 N$9193 N$9194 "Straight Waveguide" sch_x=-3 sch_y=-14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4598 N$9195 N$9196 "Straight Waveguide" sch_x=-4 sch_y=-15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4599 N$9197 N$9198 "Straight Waveguide" sch_x=0 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4600 N$9199 N$9200 "Straight Waveguide" sch_x=-1 sch_y=-12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4601 N$9201 N$9202 "Straight Waveguide" sch_x=-1 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4602 N$9203 N$9204 "Straight Waveguide" sch_x=1 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4603 N$9205 N$9206 "Straight Waveguide" sch_x=1 sch_y=-12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4604 N$9207 N$9208 "Straight Waveguide" sch_x=0 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4605 N$9209 N$9210 "Straight Waveguide" sch_x=0 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4606 N$9211 N$9212 "Straight Waveguide" sch_x=-1 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4607 N$9213 N$9214 "Straight Waveguide" sch_x=-1 sch_y=-15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4608 N$9215 N$9216 "Straight Waveguide" sch_x=1 sch_y=-15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4609 N$9217 N$9218 "Straight Waveguide" sch_x=1 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4610 N$9219 N$9220 "Straight Waveguide" sch_x=0 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4611 N$9221 N$9222 "Straight Waveguide" sch_x=4 sch_y=-12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4612 N$9223 N$9224 "Straight Waveguide" sch_x=3 sch_y=-13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4613 N$9225 N$9226 "Straight Waveguide" sch_x=3 sch_y=-14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4614 N$9227 N$9228 "Straight Waveguide" sch_x=5 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4615 N$9229 N$9230 "Straight Waveguide" sch_x=5 sch_y=-13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4616 N$9231 N$9232 "Straight Waveguide" sch_x=4 sch_y=-15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4617 N$9234 N$9233 "Straight Waveguide" sch_x=-13 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4618 N$9236 N$9235 "Straight Waveguide" sch_x=-13 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4619 N$9238 N$9237 "Straight Waveguide" sch_x=-13 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4620 N$9240 N$9239 "Straight Waveguide" sch_x=-13 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4621 N$9242 N$9241 "Straight Waveguide" sch_x=-13 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4622 N$9244 N$9243 "Straight Waveguide" sch_x=-13 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4623 N$9246 N$9245 "Straight Waveguide" sch_x=-11 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4624 N$9248 N$9247 "Straight Waveguide" sch_x=-11 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4625 N$9250 N$9249 "Straight Waveguide" sch_x=-11 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4626 N$9252 N$9251 "Straight Waveguide" sch_x=-11 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4627 N$9254 N$9253 "Straight Waveguide" sch_x=-9 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4628 N$9256 N$9255 "Straight Waveguide" sch_x=-9 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4629 N$9257 N$9258 "Straight Waveguide" sch_x=-9 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4630 N$9259 N$9260 "Straight Waveguide" sch_x=-8 sch_y=-10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4631 N$9261 N$9262 "Straight Waveguide" sch_x=-7 sch_y=-11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4632 N$9263 N$9264 "Straight Waveguide" sch_x=-7 sch_y=-12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4633 N$9265 N$9266 "Straight Waveguide" sch_x=-8 sch_y=-13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4634 N$9267 N$9268 "Straight Waveguide" sch_x=-9 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4635 N$9269 N$9270 "Straight Waveguide" sch_x=-10 sch_y=-9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4636 N$9271 N$9272 "Straight Waveguide" sch_x=-10 sch_y=-14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4637 N$9273 N$9274 "Straight Waveguide" sch_x=13 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4638 N$9275 N$9276 "Straight Waveguide" sch_x=13 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4639 N$9277 N$9278 "Straight Waveguide" sch_x=13 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4640 N$9279 N$9280 "Straight Waveguide" sch_x=13 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4641 N$9281 N$9282 "Straight Waveguide" sch_x=13 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4642 N$9283 N$9284 "Straight Waveguide" sch_x=13 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4643 N$9285 N$9286 "Straight Waveguide" sch_x=11 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4644 N$9287 N$9288 "Straight Waveguide" sch_x=11 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4645 N$9289 N$9290 "Straight Waveguide" sch_x=11 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4646 N$9291 N$9292 "Straight Waveguide" sch_x=11 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4647 N$9293 N$9294 "Straight Waveguide" sch_x=9 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4648 N$9295 N$9296 "Straight Waveguide" sch_x=9 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4649 N$9298 N$9297 "Straight Waveguide" sch_x=9 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4650 N$9300 N$9299 "Straight Waveguide" sch_x=8 sch_y=-10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4651 N$9302 N$9301 "Straight Waveguide" sch_x=7 sch_y=-11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4652 N$9304 N$9303 "Straight Waveguide" sch_x=7 sch_y=-12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4653 N$9306 N$9305 "Straight Waveguide" sch_x=8 sch_y=-13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4654 N$9308 N$9307 "Straight Waveguide" sch_x=9 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4655 N$9310 N$9309 "Straight Waveguide" sch_x=10 sch_y=-9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4656 N$9312 N$9311 "Straight Waveguide" sch_x=10 sch_y=-14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4657 N$9314 N$9313 "Straight Waveguide" sch_x=-29 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4658 N$9316 N$9315 "Straight Waveguide" sch_x=-29 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4659 N$9318 N$9317 "Straight Waveguide" sch_x=-29 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4660 N$9320 N$9319 "Straight Waveguide" sch_x=-29 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4661 N$9322 N$9321 "Straight Waveguide" sch_x=-29 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4662 N$9324 N$9323 "Straight Waveguide" sch_x=-29 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4663 N$9326 N$9325 "Straight Waveguide" sch_x=-29 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4664 N$9328 N$9327 "Straight Waveguide" sch_x=-29 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4665 N$9330 N$9329 "Straight Waveguide" sch_x=-29 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4666 N$9332 N$9331 "Straight Waveguide" sch_x=-29 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4667 N$9334 N$9333 "Straight Waveguide" sch_x=-29 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4668 N$9336 N$9335 "Straight Waveguide" sch_x=-29 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4669 N$9338 N$9337 "Straight Waveguide" sch_x=-29 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4670 N$9340 N$9339 "Straight Waveguide" sch_x=-29 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4671 N$9342 N$9341 "Straight Waveguide" sch_x=-27 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4672 N$9344 N$9343 "Straight Waveguide" sch_x=-27 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4673 N$9346 N$9345 "Straight Waveguide" sch_x=-27 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4674 N$9348 N$9347 "Straight Waveguide" sch_x=-27 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4675 N$9350 N$9349 "Straight Waveguide" sch_x=-27 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4676 N$9352 N$9351 "Straight Waveguide" sch_x=-27 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4677 N$9354 N$9353 "Straight Waveguide" sch_x=-27 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4678 N$9356 N$9355 "Straight Waveguide" sch_x=-27 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4679 N$9358 N$9357 "Straight Waveguide" sch_x=-27 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4680 N$9360 N$9359 "Straight Waveguide" sch_x=-27 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4681 N$9362 N$9361 "Straight Waveguide" sch_x=-27 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4682 N$9364 N$9363 "Straight Waveguide" sch_x=-27 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4683 N$9366 N$9365 "Straight Waveguide" sch_x=-25 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4684 N$9368 N$9367 "Straight Waveguide" sch_x=-25 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4685 N$9370 N$9369 "Straight Waveguide" sch_x=-25 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4686 N$9372 N$9371 "Straight Waveguide" sch_x=-25 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4687 N$9374 N$9373 "Straight Waveguide" sch_x=-25 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4688 N$9376 N$9375 "Straight Waveguide" sch_x=-25 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4689 N$9378 N$9377 "Straight Waveguide" sch_x=-25 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4690 N$9380 N$9379 "Straight Waveguide" sch_x=-25 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4691 N$9382 N$9381 "Straight Waveguide" sch_x=-25 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4692 N$9384 N$9383 "Straight Waveguide" sch_x=-25 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4693 N$9386 N$9385 "Straight Waveguide" sch_x=-23 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4694 N$9388 N$9387 "Straight Waveguide" sch_x=-23 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4695 N$9390 N$9389 "Straight Waveguide" sch_x=-23 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4696 N$9392 N$9391 "Straight Waveguide" sch_x=-23 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4697 N$9394 N$9393 "Straight Waveguide" sch_x=-23 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4698 N$9396 N$9395 "Straight Waveguide" sch_x=-23 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4699 N$9398 N$9397 "Straight Waveguide" sch_x=-23 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4700 N$9400 N$9399 "Straight Waveguide" sch_x=-23 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4701 N$9402 N$9401 "Straight Waveguide" sch_x=-21 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4702 N$9404 N$9403 "Straight Waveguide" sch_x=-21 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4703 N$9406 N$9405 "Straight Waveguide" sch_x=-21 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4704 N$9408 N$9407 "Straight Waveguide" sch_x=-21 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4705 N$9410 N$9409 "Straight Waveguide" sch_x=-21 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4706 N$9412 N$9411 "Straight Waveguide" sch_x=-21 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4707 N$9414 N$9413 "Straight Waveguide" sch_x=-19 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4708 N$9416 N$9415 "Straight Waveguide" sch_x=-19 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4709 N$9418 N$9417 "Straight Waveguide" sch_x=-19 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4710 N$9420 N$9419 "Straight Waveguide" sch_x=-19 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4711 N$9422 N$9421 "Straight Waveguide" sch_x=-17 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4712 N$9424 N$9423 "Straight Waveguide" sch_x=-17 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4713 N$9425 N$9426 "Straight Waveguide" sch_x=-21 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4714 N$9427 N$9428 "Straight Waveguide" sch_x=-20 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4715 N$9429 N$9430 "Straight Waveguide" sch_x=-19 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4716 N$9431 N$9432 "Straight Waveguide" sch_x=-18 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4717 N$9433 N$9434 "Straight Waveguide" sch_x=-17 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4718 N$9435 N$9436 "Straight Waveguide" sch_x=-16 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4719 N$9437 N$9438 "Straight Waveguide" sch_x=-15 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4720 N$9439 N$9440 "Straight Waveguide" sch_x=-15 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4721 N$9441 N$9442 "Straight Waveguide" sch_x=-16 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4722 N$9443 N$9444 "Straight Waveguide" sch_x=-17 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4723 N$9445 N$9446 "Straight Waveguide" sch_x=-18 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4724 N$9447 N$9448 "Straight Waveguide" sch_x=-19 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4725 N$9449 N$9450 "Straight Waveguide" sch_x=-20 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4726 N$9451 N$9452 "Straight Waveguide" sch_x=-21 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4727 N$9453 N$9454 "Straight Waveguide" sch_x=-22 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4728 N$9455 N$9456 "Straight Waveguide" sch_x=-22 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4729 N$9457 N$9458 "Straight Waveguide" sch_x=29 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4730 N$9459 N$9460 "Straight Waveguide" sch_x=29 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4731 N$9461 N$9462 "Straight Waveguide" sch_x=29 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4732 N$9463 N$9464 "Straight Waveguide" sch_x=29 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4733 N$9465 N$9466 "Straight Waveguide" sch_x=29 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4734 N$9467 N$9468 "Straight Waveguide" sch_x=29 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4735 N$9469 N$9470 "Straight Waveguide" sch_x=29 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4736 N$9471 N$9472 "Straight Waveguide" sch_x=29 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4737 N$9473 N$9474 "Straight Waveguide" sch_x=29 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4738 N$9475 N$9476 "Straight Waveguide" sch_x=29 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4739 N$9477 N$9478 "Straight Waveguide" sch_x=29 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4740 N$9479 N$9480 "Straight Waveguide" sch_x=29 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4741 N$9481 N$9482 "Straight Waveguide" sch_x=29 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4742 N$9483 N$9484 "Straight Waveguide" sch_x=29 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4743 N$9485 N$9486 "Straight Waveguide" sch_x=27 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4744 N$9487 N$9488 "Straight Waveguide" sch_x=27 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4745 N$9489 N$9490 "Straight Waveguide" sch_x=27 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4746 N$9491 N$9492 "Straight Waveguide" sch_x=27 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4747 N$9493 N$9494 "Straight Waveguide" sch_x=27 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4748 N$9495 N$9496 "Straight Waveguide" sch_x=27 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4749 N$9497 N$9498 "Straight Waveguide" sch_x=27 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4750 N$9499 N$9500 "Straight Waveguide" sch_x=27 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4751 N$9501 N$9502 "Straight Waveguide" sch_x=27 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4752 N$9503 N$9504 "Straight Waveguide" sch_x=27 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4753 N$9505 N$9506 "Straight Waveguide" sch_x=27 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4754 N$9507 N$9508 "Straight Waveguide" sch_x=27 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4755 N$9509 N$9510 "Straight Waveguide" sch_x=25 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4756 N$9511 N$9512 "Straight Waveguide" sch_x=25 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4757 N$9513 N$9514 "Straight Waveguide" sch_x=25 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4758 N$9515 N$9516 "Straight Waveguide" sch_x=25 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4759 N$9517 N$9518 "Straight Waveguide" sch_x=25 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4760 N$9519 N$9520 "Straight Waveguide" sch_x=25 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4761 N$9521 N$9522 "Straight Waveguide" sch_x=25 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4762 N$9523 N$9524 "Straight Waveguide" sch_x=25 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4763 N$9525 N$9526 "Straight Waveguide" sch_x=25 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4764 N$9527 N$9528 "Straight Waveguide" sch_x=25 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4765 N$9529 N$9530 "Straight Waveguide" sch_x=23 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4766 N$9531 N$9532 "Straight Waveguide" sch_x=23 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4767 N$9533 N$9534 "Straight Waveguide" sch_x=23 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4768 N$9535 N$9536 "Straight Waveguide" sch_x=23 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4769 N$9537 N$9538 "Straight Waveguide" sch_x=23 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4770 N$9539 N$9540 "Straight Waveguide" sch_x=23 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4771 N$9541 N$9542 "Straight Waveguide" sch_x=23 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4772 N$9543 N$9544 "Straight Waveguide" sch_x=23 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4773 N$9545 N$9546 "Straight Waveguide" sch_x=21 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4774 N$9547 N$9548 "Straight Waveguide" sch_x=21 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4775 N$9549 N$9550 "Straight Waveguide" sch_x=21 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4776 N$9551 N$9552 "Straight Waveguide" sch_x=21 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4777 N$9553 N$9554 "Straight Waveguide" sch_x=21 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4778 N$9555 N$9556 "Straight Waveguide" sch_x=21 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4779 N$9557 N$9558 "Straight Waveguide" sch_x=19 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4780 N$9559 N$9560 "Straight Waveguide" sch_x=19 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4781 N$9561 N$9562 "Straight Waveguide" sch_x=19 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4782 N$9563 N$9564 "Straight Waveguide" sch_x=19 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4783 N$9565 N$9566 "Straight Waveguide" sch_x=17 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4784 N$9567 N$9568 "Straight Waveguide" sch_x=17 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4785 N$9570 N$9569 "Straight Waveguide" sch_x=21 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4786 N$9572 N$9571 "Straight Waveguide" sch_x=20 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4787 N$9574 N$9573 "Straight Waveguide" sch_x=19 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4788 N$9576 N$9575 "Straight Waveguide" sch_x=18 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4789 N$9578 N$9577 "Straight Waveguide" sch_x=17 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4790 N$9580 N$9579 "Straight Waveguide" sch_x=16 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4791 N$9582 N$9581 "Straight Waveguide" sch_x=15 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4792 N$9584 N$9583 "Straight Waveguide" sch_x=15 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4793 N$9586 N$9585 "Straight Waveguide" sch_x=16 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4794 N$9588 N$9587 "Straight Waveguide" sch_x=17 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4795 N$9590 N$9589 "Straight Waveguide" sch_x=18 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4796 N$9592 N$9591 "Straight Waveguide" sch_x=19 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4797 N$9594 N$9593 "Straight Waveguide" sch_x=20 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4798 N$9596 N$9595 "Straight Waveguide" sch_x=21 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4799 N$9598 N$9597 "Straight Waveguide" sch_x=22 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4800 N$9600 N$9599 "Straight Waveguide" sch_x=22 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4801 N$9601 N$9602 "Straight Waveguide" sch_x=-4 sch_y=-16.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4802 N$9603 N$9604 "Straight Waveguide" sch_x=-5 sch_y=-17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4803 N$9605 N$9606 "Straight Waveguide" sch_x=-5 sch_y=-18.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4804 N$9607 N$9608 "Straight Waveguide" sch_x=-3 sch_y=-17.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4805 N$9609 N$9610 "Straight Waveguide" sch_x=-3 sch_y=-18.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4806 N$9611 N$9612 "Straight Waveguide" sch_x=-4 sch_y=-19.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4807 N$9613 N$9614 "Straight Waveguide" sch_x=0 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4808 N$9615 N$9616 "Straight Waveguide" sch_x=-1 sch_y=-16.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4809 N$9617 N$9618 "Straight Waveguide" sch_x=-1 sch_y=-17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4810 N$9619 N$9620 "Straight Waveguide" sch_x=1 sch_y=-17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4811 N$9621 N$9622 "Straight Waveguide" sch_x=1 sch_y=-16.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4812 N$9623 N$9624 "Straight Waveguide" sch_x=0 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4813 N$9625 N$9626 "Straight Waveguide" sch_x=0 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4814 N$9627 N$9628 "Straight Waveguide" sch_x=-1 sch_y=-18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4815 N$9629 N$9630 "Straight Waveguide" sch_x=-1 sch_y=-19.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4816 N$9631 N$9632 "Straight Waveguide" sch_x=1 sch_y=-19.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4817 N$9633 N$9634 "Straight Waveguide" sch_x=1 sch_y=-18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4818 N$9635 N$9636 "Straight Waveguide" sch_x=0 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4819 N$9637 N$9638 "Straight Waveguide" sch_x=4 sch_y=-16.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4820 N$9639 N$9640 "Straight Waveguide" sch_x=3 sch_y=-17.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4821 N$9641 N$9642 "Straight Waveguide" sch_x=3 sch_y=-18.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4822 N$9643 N$9644 "Straight Waveguide" sch_x=5 sch_y=-18.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4823 N$9645 N$9646 "Straight Waveguide" sch_x=5 sch_y=-17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4824 N$9647 N$9648 "Straight Waveguide" sch_x=4 sch_y=-19.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4825 N$9649 N$9650 "Straight Waveguide" sch_x=-4 sch_y=-20.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4826 N$9651 N$9652 "Straight Waveguide" sch_x=-5 sch_y=-21.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4827 N$9653 N$9654 "Straight Waveguide" sch_x=-5 sch_y=-22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4828 N$9655 N$9656 "Straight Waveguide" sch_x=-3 sch_y=-21.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4829 N$9657 N$9658 "Straight Waveguide" sch_x=-3 sch_y=-22.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4830 N$9659 N$9660 "Straight Waveguide" sch_x=-4 sch_y=-23.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4831 N$9661 N$9662 "Straight Waveguide" sch_x=0 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4832 N$9663 N$9664 "Straight Waveguide" sch_x=-1 sch_y=-20.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4833 N$9665 N$9666 "Straight Waveguide" sch_x=-1 sch_y=-21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4834 N$9667 N$9668 "Straight Waveguide" sch_x=1 sch_y=-21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4835 N$9669 N$9670 "Straight Waveguide" sch_x=1 sch_y=-20.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4836 N$9671 N$9672 "Straight Waveguide" sch_x=0 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4837 N$9673 N$9674 "Straight Waveguide" sch_x=0 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4838 N$9675 N$9676 "Straight Waveguide" sch_x=-1 sch_y=-22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4839 N$9677 N$9678 "Straight Waveguide" sch_x=-1 sch_y=-23.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4840 N$9679 N$9680 "Straight Waveguide" sch_x=1 sch_y=-23.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4841 N$9681 N$9682 "Straight Waveguide" sch_x=1 sch_y=-22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4842 N$9683 N$9684 "Straight Waveguide" sch_x=0 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4843 N$9685 N$9686 "Straight Waveguide" sch_x=4 sch_y=-20.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4844 N$9687 N$9688 "Straight Waveguide" sch_x=3 sch_y=-21.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4845 N$9689 N$9690 "Straight Waveguide" sch_x=3 sch_y=-22.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4846 N$9691 N$9692 "Straight Waveguide" sch_x=5 sch_y=-22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4847 N$9693 N$9694 "Straight Waveguide" sch_x=5 sch_y=-21.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4848 N$9695 N$9696 "Straight Waveguide" sch_x=4 sch_y=-23.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4849 N$9698 N$9697 "Straight Waveguide" sch_x=-13 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4850 N$9700 N$9699 "Straight Waveguide" sch_x=-13 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4851 N$9702 N$9701 "Straight Waveguide" sch_x=-13 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4852 N$9704 N$9703 "Straight Waveguide" sch_x=-13 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4853 N$9706 N$9705 "Straight Waveguide" sch_x=-13 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4854 N$9708 N$9707 "Straight Waveguide" sch_x=-13 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4855 N$9710 N$9709 "Straight Waveguide" sch_x=-11 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4856 N$9712 N$9711 "Straight Waveguide" sch_x=-11 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4857 N$9714 N$9713 "Straight Waveguide" sch_x=-11 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4858 N$9716 N$9715 "Straight Waveguide" sch_x=-11 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4859 N$9718 N$9717 "Straight Waveguide" sch_x=-9 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4860 N$9720 N$9719 "Straight Waveguide" sch_x=-9 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4861 N$9721 N$9722 "Straight Waveguide" sch_x=-9 sch_y=-17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4862 N$9723 N$9724 "Straight Waveguide" sch_x=-8 sch_y=-18.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4863 N$9725 N$9726 "Straight Waveguide" sch_x=-7 sch_y=-19.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4864 N$9727 N$9728 "Straight Waveguide" sch_x=-7 sch_y=-20.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4865 N$9729 N$9730 "Straight Waveguide" sch_x=-8 sch_y=-21.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4866 N$9731 N$9732 "Straight Waveguide" sch_x=-9 sch_y=-22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4867 N$9733 N$9734 "Straight Waveguide" sch_x=-10 sch_y=-17.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4868 N$9735 N$9736 "Straight Waveguide" sch_x=-10 sch_y=-22.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4869 N$9737 N$9738 "Straight Waveguide" sch_x=13 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4870 N$9739 N$9740 "Straight Waveguide" sch_x=13 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4871 N$9741 N$9742 "Straight Waveguide" sch_x=13 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4872 N$9743 N$9744 "Straight Waveguide" sch_x=13 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4873 N$9745 N$9746 "Straight Waveguide" sch_x=13 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4874 N$9747 N$9748 "Straight Waveguide" sch_x=13 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4875 N$9749 N$9750 "Straight Waveguide" sch_x=11 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4876 N$9751 N$9752 "Straight Waveguide" sch_x=11 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4877 N$9753 N$9754 "Straight Waveguide" sch_x=11 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4878 N$9755 N$9756 "Straight Waveguide" sch_x=11 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4879 N$9757 N$9758 "Straight Waveguide" sch_x=9 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4880 N$9759 N$9760 "Straight Waveguide" sch_x=9 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4881 N$9762 N$9761 "Straight Waveguide" sch_x=9 sch_y=-17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4882 N$9764 N$9763 "Straight Waveguide" sch_x=8 sch_y=-18.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4883 N$9766 N$9765 "Straight Waveguide" sch_x=7 sch_y=-19.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4884 N$9768 N$9767 "Straight Waveguide" sch_x=7 sch_y=-20.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4885 N$9770 N$9769 "Straight Waveguide" sch_x=8 sch_y=-21.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4886 N$9772 N$9771 "Straight Waveguide" sch_x=9 sch_y=-22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4887 N$9774 N$9773 "Straight Waveguide" sch_x=10 sch_y=-17.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4888 N$9776 N$9775 "Straight Waveguide" sch_x=10 sch_y=-22.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4889 N$9777 N$9778 "Straight Waveguide" sch_x=-4 sch_y=-24.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4890 N$9779 N$9780 "Straight Waveguide" sch_x=-5 sch_y=-25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4891 N$9781 N$9782 "Straight Waveguide" sch_x=-5 sch_y=-26.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4892 N$9783 N$9784 "Straight Waveguide" sch_x=-3 sch_y=-25.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4893 N$9785 N$9786 "Straight Waveguide" sch_x=-3 sch_y=-26.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4894 N$9787 N$9788 "Straight Waveguide" sch_x=-4 sch_y=-27.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4895 N$9789 N$9790 "Straight Waveguide" sch_x=0 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4896 N$9791 N$9792 "Straight Waveguide" sch_x=-1 sch_y=-24.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4897 N$9793 N$9794 "Straight Waveguide" sch_x=-1 sch_y=-25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4898 N$9795 N$9796 "Straight Waveguide" sch_x=1 sch_y=-25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4899 N$9797 N$9798 "Straight Waveguide" sch_x=1 sch_y=-24.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4900 N$9799 N$9800 "Straight Waveguide" sch_x=0 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4901 N$9801 N$9802 "Straight Waveguide" sch_x=0 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4902 N$9803 N$9804 "Straight Waveguide" sch_x=-1 sch_y=-26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4903 N$9805 N$9806 "Straight Waveguide" sch_x=-1 sch_y=-27.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4904 N$9807 N$9808 "Straight Waveguide" sch_x=1 sch_y=-27.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4905 N$9809 N$9810 "Straight Waveguide" sch_x=1 sch_y=-26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4906 N$9811 N$9812 "Straight Waveguide" sch_x=0 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4907 N$9813 N$9814 "Straight Waveguide" sch_x=4 sch_y=-24.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4908 N$9815 N$9816 "Straight Waveguide" sch_x=3 sch_y=-25.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4909 N$9817 N$9818 "Straight Waveguide" sch_x=3 sch_y=-26.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4910 N$9819 N$9820 "Straight Waveguide" sch_x=5 sch_y=-26.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4911 N$9821 N$9822 "Straight Waveguide" sch_x=5 sch_y=-25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4912 N$9823 N$9824 "Straight Waveguide" sch_x=4 sch_y=-27.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4913 N$9825 N$9826 "Straight Waveguide" sch_x=-4 sch_y=-28.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4914 N$9827 N$9828 "Straight Waveguide" sch_x=-5 sch_y=-29.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4915 N$9829 N$9830 "Straight Waveguide" sch_x=-5 sch_y=-30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4916 N$9831 N$9832 "Straight Waveguide" sch_x=-3 sch_y=-29.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4917 N$9833 N$9834 "Straight Waveguide" sch_x=-3 sch_y=-30.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4918 N$9835 N$9836 "Straight Waveguide" sch_x=-4 sch_y=-31.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4919 N$9837 N$9838 "Straight Waveguide" sch_x=0 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4920 N$9839 N$9840 "Straight Waveguide" sch_x=-1 sch_y=-28.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4921 N$9841 N$9842 "Straight Waveguide" sch_x=-1 sch_y=-29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4922 N$9843 N$9844 "Straight Waveguide" sch_x=1 sch_y=-29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4923 N$9845 N$9846 "Straight Waveguide" sch_x=1 sch_y=-28.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4924 N$9847 N$9848 "Straight Waveguide" sch_x=0 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4925 N$9849 N$9850 "Straight Waveguide" sch_x=0 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4926 N$9851 N$9852 "Straight Waveguide" sch_x=-1 sch_y=-30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4927 N$9853 N$9854 "Straight Waveguide" sch_x=-1 sch_y=-31.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4928 N$9855 N$9856 "Straight Waveguide" sch_x=1 sch_y=-31.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4929 N$9857 N$9858 "Straight Waveguide" sch_x=1 sch_y=-30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4930 N$9859 N$9860 "Straight Waveguide" sch_x=0 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4931 N$9861 N$9862 "Straight Waveguide" sch_x=4 sch_y=-28.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4932 N$9863 N$9864 "Straight Waveguide" sch_x=3 sch_y=-29.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4933 N$9865 N$9866 "Straight Waveguide" sch_x=3 sch_y=-30.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4934 N$9867 N$9868 "Straight Waveguide" sch_x=5 sch_y=-30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4935 N$9869 N$9870 "Straight Waveguide" sch_x=5 sch_y=-29.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4936 N$9871 N$9872 "Straight Waveguide" sch_x=4 sch_y=-31.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4937 N$9874 N$9873 "Straight Waveguide" sch_x=-13 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4938 N$9876 N$9875 "Straight Waveguide" sch_x=-13 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4939 N$9878 N$9877 "Straight Waveguide" sch_x=-13 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4940 N$9880 N$9879 "Straight Waveguide" sch_x=-13 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4941 N$9882 N$9881 "Straight Waveguide" sch_x=-13 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4942 N$9884 N$9883 "Straight Waveguide" sch_x=-13 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4943 N$9886 N$9885 "Straight Waveguide" sch_x=-11 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4944 N$9888 N$9887 "Straight Waveguide" sch_x=-11 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4945 N$9890 N$9889 "Straight Waveguide" sch_x=-11 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4946 N$9892 N$9891 "Straight Waveguide" sch_x=-11 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4947 N$9894 N$9893 "Straight Waveguide" sch_x=-9 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4948 N$9896 N$9895 "Straight Waveguide" sch_x=-9 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4949 N$9897 N$9898 "Straight Waveguide" sch_x=-9 sch_y=-25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4950 N$9899 N$9900 "Straight Waveguide" sch_x=-8 sch_y=-26.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4951 N$9901 N$9902 "Straight Waveguide" sch_x=-7 sch_y=-27.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4952 N$9903 N$9904 "Straight Waveguide" sch_x=-7 sch_y=-28.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4953 N$9905 N$9906 "Straight Waveguide" sch_x=-8 sch_y=-29.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4954 N$9907 N$9908 "Straight Waveguide" sch_x=-9 sch_y=-30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4955 N$9909 N$9910 "Straight Waveguide" sch_x=-10 sch_y=-25.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4956 N$9911 N$9912 "Straight Waveguide" sch_x=-10 sch_y=-30.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4957 N$9913 N$9914 "Straight Waveguide" sch_x=13 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4958 N$9915 N$9916 "Straight Waveguide" sch_x=13 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4959 N$9917 N$9918 "Straight Waveguide" sch_x=13 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4960 N$9919 N$9920 "Straight Waveguide" sch_x=13 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4961 N$9921 N$9922 "Straight Waveguide" sch_x=13 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4962 N$9923 N$9924 "Straight Waveguide" sch_x=13 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4963 N$9925 N$9926 "Straight Waveguide" sch_x=11 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4964 N$9927 N$9928 "Straight Waveguide" sch_x=11 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4965 N$9929 N$9930 "Straight Waveguide" sch_x=11 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4966 N$9931 N$9932 "Straight Waveguide" sch_x=11 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4967 N$9933 N$9934 "Straight Waveguide" sch_x=9 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4968 N$9935 N$9936 "Straight Waveguide" sch_x=9 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4969 N$9938 N$9937 "Straight Waveguide" sch_x=9 sch_y=-25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4970 N$9940 N$9939 "Straight Waveguide" sch_x=8 sch_y=-26.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4971 N$9942 N$9941 "Straight Waveguide" sch_x=7 sch_y=-27.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4972 N$9944 N$9943 "Straight Waveguide" sch_x=7 sch_y=-28.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4973 N$9946 N$9945 "Straight Waveguide" sch_x=8 sch_y=-29.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4974 N$9948 N$9947 "Straight Waveguide" sch_x=9 sch_y=-30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4975 N$9950 N$9949 "Straight Waveguide" sch_x=10 sch_y=-25.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4976 N$9952 N$9951 "Straight Waveguide" sch_x=10 sch_y=-30.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4977 N$9954 N$9953 "Straight Waveguide" sch_x=-29 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4978 N$9956 N$9955 "Straight Waveguide" sch_x=-29 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4979 N$9958 N$9957 "Straight Waveguide" sch_x=-29 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4980 N$9960 N$9959 "Straight Waveguide" sch_x=-29 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4981 N$9962 N$9961 "Straight Waveguide" sch_x=-29 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4982 N$9964 N$9963 "Straight Waveguide" sch_x=-29 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4983 N$9966 N$9965 "Straight Waveguide" sch_x=-29 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4984 N$9968 N$9967 "Straight Waveguide" sch_x=-29 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4985 N$9970 N$9969 "Straight Waveguide" sch_x=-29 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4986 N$9972 N$9971 "Straight Waveguide" sch_x=-29 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4987 N$9974 N$9973 "Straight Waveguide" sch_x=-29 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4988 N$9976 N$9975 "Straight Waveguide" sch_x=-29 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4989 N$9978 N$9977 "Straight Waveguide" sch_x=-29 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4990 N$9980 N$9979 "Straight Waveguide" sch_x=-29 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4991 N$9982 N$9981 "Straight Waveguide" sch_x=-27 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4992 N$9984 N$9983 "Straight Waveguide" sch_x=-27 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4993 N$9986 N$9985 "Straight Waveguide" sch_x=-27 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4994 N$9988 N$9987 "Straight Waveguide" sch_x=-27 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4995 N$9990 N$9989 "Straight Waveguide" sch_x=-27 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4996 N$9992 N$9991 "Straight Waveguide" sch_x=-27 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4997 N$9994 N$9993 "Straight Waveguide" sch_x=-27 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4998 N$9996 N$9995 "Straight Waveguide" sch_x=-27 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4999 N$9998 N$9997 "Straight Waveguide" sch_x=-27 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5000 N$10000 N$9999 "Straight Waveguide" sch_x=-27 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5001 N$10002 N$10001 "Straight Waveguide" sch_x=-27 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5002 N$10004 N$10003 "Straight Waveguide" sch_x=-27 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5003 N$10006 N$10005 "Straight Waveguide" sch_x=-25 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5004 N$10008 N$10007 "Straight Waveguide" sch_x=-25 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5005 N$10010 N$10009 "Straight Waveguide" sch_x=-25 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5006 N$10012 N$10011 "Straight Waveguide" sch_x=-25 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5007 N$10014 N$10013 "Straight Waveguide" sch_x=-25 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5008 N$10016 N$10015 "Straight Waveguide" sch_x=-25 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5009 N$10018 N$10017 "Straight Waveguide" sch_x=-25 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5010 N$10020 N$10019 "Straight Waveguide" sch_x=-25 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5011 N$10022 N$10021 "Straight Waveguide" sch_x=-25 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5012 N$10024 N$10023 "Straight Waveguide" sch_x=-25 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5013 N$10026 N$10025 "Straight Waveguide" sch_x=-23 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5014 N$10028 N$10027 "Straight Waveguide" sch_x=-23 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5015 N$10030 N$10029 "Straight Waveguide" sch_x=-23 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5016 N$10032 N$10031 "Straight Waveguide" sch_x=-23 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5017 N$10034 N$10033 "Straight Waveguide" sch_x=-23 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5018 N$10036 N$10035 "Straight Waveguide" sch_x=-23 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5019 N$10038 N$10037 "Straight Waveguide" sch_x=-23 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5020 N$10040 N$10039 "Straight Waveguide" sch_x=-23 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5021 N$10042 N$10041 "Straight Waveguide" sch_x=-21 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5022 N$10044 N$10043 "Straight Waveguide" sch_x=-21 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5023 N$10046 N$10045 "Straight Waveguide" sch_x=-21 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5024 N$10048 N$10047 "Straight Waveguide" sch_x=-21 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5025 N$10050 N$10049 "Straight Waveguide" sch_x=-21 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5026 N$10052 N$10051 "Straight Waveguide" sch_x=-21 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5027 N$10054 N$10053 "Straight Waveguide" sch_x=-19 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5028 N$10056 N$10055 "Straight Waveguide" sch_x=-19 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5029 N$10058 N$10057 "Straight Waveguide" sch_x=-19 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5030 N$10060 N$10059 "Straight Waveguide" sch_x=-19 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5031 N$10062 N$10061 "Straight Waveguide" sch_x=-17 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5032 N$10064 N$10063 "Straight Waveguide" sch_x=-17 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5033 N$10065 N$10066 "Straight Waveguide" sch_x=-21 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5034 N$10067 N$10068 "Straight Waveguide" sch_x=-20 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5035 N$10069 N$10070 "Straight Waveguide" sch_x=-19 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5036 N$10071 N$10072 "Straight Waveguide" sch_x=-18 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5037 N$10073 N$10074 "Straight Waveguide" sch_x=-17 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5038 N$10075 N$10076 "Straight Waveguide" sch_x=-16 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5039 N$10077 N$10078 "Straight Waveguide" sch_x=-15 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5040 N$10079 N$10080 "Straight Waveguide" sch_x=-15 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5041 N$10081 N$10082 "Straight Waveguide" sch_x=-16 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5042 N$10083 N$10084 "Straight Waveguide" sch_x=-17 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5043 N$10085 N$10086 "Straight Waveguide" sch_x=-18 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5044 N$10087 N$10088 "Straight Waveguide" sch_x=-19 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5045 N$10089 N$10090 "Straight Waveguide" sch_x=-20 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5046 N$10091 N$10092 "Straight Waveguide" sch_x=-21 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5047 N$10093 N$10094 "Straight Waveguide" sch_x=-22 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5048 N$10095 N$10096 "Straight Waveguide" sch_x=-22 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5049 N$10097 N$10098 "Straight Waveguide" sch_x=29 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5050 N$10099 N$10100 "Straight Waveguide" sch_x=29 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5051 N$10101 N$10102 "Straight Waveguide" sch_x=29 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5052 N$10103 N$10104 "Straight Waveguide" sch_x=29 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5053 N$10105 N$10106 "Straight Waveguide" sch_x=29 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5054 N$10107 N$10108 "Straight Waveguide" sch_x=29 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5055 N$10109 N$10110 "Straight Waveguide" sch_x=29 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5056 N$10111 N$10112 "Straight Waveguide" sch_x=29 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5057 N$10113 N$10114 "Straight Waveguide" sch_x=29 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5058 N$10115 N$10116 "Straight Waveguide" sch_x=29 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5059 N$10117 N$10118 "Straight Waveguide" sch_x=29 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5060 N$10119 N$10120 "Straight Waveguide" sch_x=29 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5061 N$10121 N$10122 "Straight Waveguide" sch_x=29 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5062 N$10123 N$10124 "Straight Waveguide" sch_x=29 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5063 N$10125 N$10126 "Straight Waveguide" sch_x=27 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5064 N$10127 N$10128 "Straight Waveguide" sch_x=27 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5065 N$10129 N$10130 "Straight Waveguide" sch_x=27 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5066 N$10131 N$10132 "Straight Waveguide" sch_x=27 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5067 N$10133 N$10134 "Straight Waveguide" sch_x=27 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5068 N$10135 N$10136 "Straight Waveguide" sch_x=27 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5069 N$10137 N$10138 "Straight Waveguide" sch_x=27 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5070 N$10139 N$10140 "Straight Waveguide" sch_x=27 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5071 N$10141 N$10142 "Straight Waveguide" sch_x=27 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5072 N$10143 N$10144 "Straight Waveguide" sch_x=27 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5073 N$10145 N$10146 "Straight Waveguide" sch_x=27 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5074 N$10147 N$10148 "Straight Waveguide" sch_x=27 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5075 N$10149 N$10150 "Straight Waveguide" sch_x=25 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5076 N$10151 N$10152 "Straight Waveguide" sch_x=25 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5077 N$10153 N$10154 "Straight Waveguide" sch_x=25 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5078 N$10155 N$10156 "Straight Waveguide" sch_x=25 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5079 N$10157 N$10158 "Straight Waveguide" sch_x=25 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5080 N$10159 N$10160 "Straight Waveguide" sch_x=25 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5081 N$10161 N$10162 "Straight Waveguide" sch_x=25 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5082 N$10163 N$10164 "Straight Waveguide" sch_x=25 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5083 N$10165 N$10166 "Straight Waveguide" sch_x=25 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5084 N$10167 N$10168 "Straight Waveguide" sch_x=25 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5085 N$10169 N$10170 "Straight Waveguide" sch_x=23 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5086 N$10171 N$10172 "Straight Waveguide" sch_x=23 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5087 N$10173 N$10174 "Straight Waveguide" sch_x=23 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5088 N$10175 N$10176 "Straight Waveguide" sch_x=23 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5089 N$10177 N$10178 "Straight Waveguide" sch_x=23 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5090 N$10179 N$10180 "Straight Waveguide" sch_x=23 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5091 N$10181 N$10182 "Straight Waveguide" sch_x=23 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5092 N$10183 N$10184 "Straight Waveguide" sch_x=23 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5093 N$10185 N$10186 "Straight Waveguide" sch_x=21 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5094 N$10187 N$10188 "Straight Waveguide" sch_x=21 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5095 N$10189 N$10190 "Straight Waveguide" sch_x=21 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5096 N$10191 N$10192 "Straight Waveguide" sch_x=21 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5097 N$10193 N$10194 "Straight Waveguide" sch_x=21 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5098 N$10195 N$10196 "Straight Waveguide" sch_x=21 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5099 N$10197 N$10198 "Straight Waveguide" sch_x=19 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5100 N$10199 N$10200 "Straight Waveguide" sch_x=19 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5101 N$10201 N$10202 "Straight Waveguide" sch_x=19 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5102 N$10203 N$10204 "Straight Waveguide" sch_x=19 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5103 N$10205 N$10206 "Straight Waveguide" sch_x=17 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5104 N$10207 N$10208 "Straight Waveguide" sch_x=17 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5105 N$10210 N$10209 "Straight Waveguide" sch_x=21 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5106 N$10212 N$10211 "Straight Waveguide" sch_x=20 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5107 N$10214 N$10213 "Straight Waveguide" sch_x=19 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5108 N$10216 N$10215 "Straight Waveguide" sch_x=18 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5109 N$10218 N$10217 "Straight Waveguide" sch_x=17 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5110 N$10220 N$10219 "Straight Waveguide" sch_x=16 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5111 N$10222 N$10221 "Straight Waveguide" sch_x=15 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5112 N$10224 N$10223 "Straight Waveguide" sch_x=15 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5113 N$10226 N$10225 "Straight Waveguide" sch_x=16 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5114 N$10228 N$10227 "Straight Waveguide" sch_x=17 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5115 N$10230 N$10229 "Straight Waveguide" sch_x=18 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5116 N$10232 N$10231 "Straight Waveguide" sch_x=19 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5117 N$10234 N$10233 "Straight Waveguide" sch_x=20 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5118 N$10236 N$10235 "Straight Waveguide" sch_x=21 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5119 N$10238 N$10237 "Straight Waveguide" sch_x=22 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5120 N$10240 N$10239 "Straight Waveguide" sch_x=22 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5121 N$10242 N$10241 "Straight Waveguide" sch_x=-61 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5122 N$10244 N$10243 "Straight Waveguide" sch_x=-61 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5123 N$10246 N$10245 "Straight Waveguide" sch_x=-61 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5124 N$10248 N$10247 "Straight Waveguide" sch_x=-61 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5125 N$10250 N$10249 "Straight Waveguide" sch_x=-61 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5126 N$10252 N$10251 "Straight Waveguide" sch_x=-61 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5127 N$10254 N$10253 "Straight Waveguide" sch_x=-61 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5128 N$10256 N$10255 "Straight Waveguide" sch_x=-61 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5129 N$10258 N$10257 "Straight Waveguide" sch_x=-61 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5130 N$10260 N$10259 "Straight Waveguide" sch_x=-61 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5131 N$10262 N$10261 "Straight Waveguide" sch_x=-61 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5132 N$10264 N$10263 "Straight Waveguide" sch_x=-61 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5133 N$10266 N$10265 "Straight Waveguide" sch_x=-61 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5134 N$10268 N$10267 "Straight Waveguide" sch_x=-61 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5135 N$10270 N$10269 "Straight Waveguide" sch_x=-61 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5136 N$10272 N$10271 "Straight Waveguide" sch_x=-61 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5137 N$10274 N$10273 "Straight Waveguide" sch_x=-61 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5138 N$10276 N$10275 "Straight Waveguide" sch_x=-61 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5139 N$10278 N$10277 "Straight Waveguide" sch_x=-61 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5140 N$10280 N$10279 "Straight Waveguide" sch_x=-61 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5141 N$10282 N$10281 "Straight Waveguide" sch_x=-61 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5142 N$10284 N$10283 "Straight Waveguide" sch_x=-61 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5143 N$10286 N$10285 "Straight Waveguide" sch_x=-61 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5144 N$10288 N$10287 "Straight Waveguide" sch_x=-61 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5145 N$10290 N$10289 "Straight Waveguide" sch_x=-61 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5146 N$10292 N$10291 "Straight Waveguide" sch_x=-61 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5147 N$10294 N$10293 "Straight Waveguide" sch_x=-61 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5148 N$10296 N$10295 "Straight Waveguide" sch_x=-61 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5149 N$10298 N$10297 "Straight Waveguide" sch_x=-61 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5150 N$10300 N$10299 "Straight Waveguide" sch_x=-61 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5151 N$10302 N$10301 "Straight Waveguide" sch_x=-59 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5152 N$10304 N$10303 "Straight Waveguide" sch_x=-59 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5153 N$10306 N$10305 "Straight Waveguide" sch_x=-59 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5154 N$10308 N$10307 "Straight Waveguide" sch_x=-59 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5155 N$10310 N$10309 "Straight Waveguide" sch_x=-59 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5156 N$10312 N$10311 "Straight Waveguide" sch_x=-59 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5157 N$10314 N$10313 "Straight Waveguide" sch_x=-59 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5158 N$10316 N$10315 "Straight Waveguide" sch_x=-59 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5159 N$10318 N$10317 "Straight Waveguide" sch_x=-59 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5160 N$10320 N$10319 "Straight Waveguide" sch_x=-59 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5161 N$10322 N$10321 "Straight Waveguide" sch_x=-59 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5162 N$10324 N$10323 "Straight Waveguide" sch_x=-59 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5163 N$10326 N$10325 "Straight Waveguide" sch_x=-59 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5164 N$10328 N$10327 "Straight Waveguide" sch_x=-59 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5165 N$10330 N$10329 "Straight Waveguide" sch_x=-59 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5166 N$10332 N$10331 "Straight Waveguide" sch_x=-59 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5167 N$10334 N$10333 "Straight Waveguide" sch_x=-59 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5168 N$10336 N$10335 "Straight Waveguide" sch_x=-59 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5169 N$10338 N$10337 "Straight Waveguide" sch_x=-59 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5170 N$10340 N$10339 "Straight Waveguide" sch_x=-59 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5171 N$10342 N$10341 "Straight Waveguide" sch_x=-59 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5172 N$10344 N$10343 "Straight Waveguide" sch_x=-59 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5173 N$10346 N$10345 "Straight Waveguide" sch_x=-59 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5174 N$10348 N$10347 "Straight Waveguide" sch_x=-59 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5175 N$10350 N$10349 "Straight Waveguide" sch_x=-59 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5176 N$10352 N$10351 "Straight Waveguide" sch_x=-59 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5177 N$10354 N$10353 "Straight Waveguide" sch_x=-59 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5178 N$10356 N$10355 "Straight Waveguide" sch_x=-59 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5179 N$10358 N$10357 "Straight Waveguide" sch_x=-57 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5180 N$10360 N$10359 "Straight Waveguide" sch_x=-57 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5181 N$10362 N$10361 "Straight Waveguide" sch_x=-57 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5182 N$10364 N$10363 "Straight Waveguide" sch_x=-57 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5183 N$10366 N$10365 "Straight Waveguide" sch_x=-57 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5184 N$10368 N$10367 "Straight Waveguide" sch_x=-57 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5185 N$10370 N$10369 "Straight Waveguide" sch_x=-57 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5186 N$10372 N$10371 "Straight Waveguide" sch_x=-57 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5187 N$10374 N$10373 "Straight Waveguide" sch_x=-57 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5188 N$10376 N$10375 "Straight Waveguide" sch_x=-57 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5189 N$10378 N$10377 "Straight Waveguide" sch_x=-57 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5190 N$10380 N$10379 "Straight Waveguide" sch_x=-57 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5191 N$10382 N$10381 "Straight Waveguide" sch_x=-57 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5192 N$10384 N$10383 "Straight Waveguide" sch_x=-57 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5193 N$10386 N$10385 "Straight Waveguide" sch_x=-57 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5194 N$10388 N$10387 "Straight Waveguide" sch_x=-57 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5195 N$10390 N$10389 "Straight Waveguide" sch_x=-57 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5196 N$10392 N$10391 "Straight Waveguide" sch_x=-57 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5197 N$10394 N$10393 "Straight Waveguide" sch_x=-57 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5198 N$10396 N$10395 "Straight Waveguide" sch_x=-57 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5199 N$10398 N$10397 "Straight Waveguide" sch_x=-57 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5200 N$10400 N$10399 "Straight Waveguide" sch_x=-57 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5201 N$10402 N$10401 "Straight Waveguide" sch_x=-57 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5202 N$10404 N$10403 "Straight Waveguide" sch_x=-57 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5203 N$10406 N$10405 "Straight Waveguide" sch_x=-57 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5204 N$10408 N$10407 "Straight Waveguide" sch_x=-57 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5205 N$10410 N$10409 "Straight Waveguide" sch_x=-55 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5206 N$10412 N$10411 "Straight Waveguide" sch_x=-55 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5207 N$10414 N$10413 "Straight Waveguide" sch_x=-55 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5208 N$10416 N$10415 "Straight Waveguide" sch_x=-55 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5209 N$10418 N$10417 "Straight Waveguide" sch_x=-55 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5210 N$10420 N$10419 "Straight Waveguide" sch_x=-55 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5211 N$10422 N$10421 "Straight Waveguide" sch_x=-55 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5212 N$10424 N$10423 "Straight Waveguide" sch_x=-55 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5213 N$10426 N$10425 "Straight Waveguide" sch_x=-55 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5214 N$10428 N$10427 "Straight Waveguide" sch_x=-55 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5215 N$10430 N$10429 "Straight Waveguide" sch_x=-55 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5216 N$10432 N$10431 "Straight Waveguide" sch_x=-55 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5217 N$10434 N$10433 "Straight Waveguide" sch_x=-55 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5218 N$10436 N$10435 "Straight Waveguide" sch_x=-55 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5219 N$10438 N$10437 "Straight Waveguide" sch_x=-55 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5220 N$10440 N$10439 "Straight Waveguide" sch_x=-55 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5221 N$10442 N$10441 "Straight Waveguide" sch_x=-55 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5222 N$10444 N$10443 "Straight Waveguide" sch_x=-55 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5223 N$10446 N$10445 "Straight Waveguide" sch_x=-55 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5224 N$10448 N$10447 "Straight Waveguide" sch_x=-55 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5225 N$10450 N$10449 "Straight Waveguide" sch_x=-55 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5226 N$10452 N$10451 "Straight Waveguide" sch_x=-55 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5227 N$10454 N$10453 "Straight Waveguide" sch_x=-55 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5228 N$10456 N$10455 "Straight Waveguide" sch_x=-55 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5229 N$10458 N$10457 "Straight Waveguide" sch_x=-53 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5230 N$10460 N$10459 "Straight Waveguide" sch_x=-53 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5231 N$10462 N$10461 "Straight Waveguide" sch_x=-53 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5232 N$10464 N$10463 "Straight Waveguide" sch_x=-53 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5233 N$10466 N$10465 "Straight Waveguide" sch_x=-53 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5234 N$10468 N$10467 "Straight Waveguide" sch_x=-53 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5235 N$10470 N$10469 "Straight Waveguide" sch_x=-53 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5236 N$10472 N$10471 "Straight Waveguide" sch_x=-53 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5237 N$10474 N$10473 "Straight Waveguide" sch_x=-53 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5238 N$10476 N$10475 "Straight Waveguide" sch_x=-53 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5239 N$10478 N$10477 "Straight Waveguide" sch_x=-53 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5240 N$10480 N$10479 "Straight Waveguide" sch_x=-53 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5241 N$10482 N$10481 "Straight Waveguide" sch_x=-53 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5242 N$10484 N$10483 "Straight Waveguide" sch_x=-53 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5243 N$10486 N$10485 "Straight Waveguide" sch_x=-53 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5244 N$10488 N$10487 "Straight Waveguide" sch_x=-53 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5245 N$10490 N$10489 "Straight Waveguide" sch_x=-53 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5246 N$10492 N$10491 "Straight Waveguide" sch_x=-53 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5247 N$10494 N$10493 "Straight Waveguide" sch_x=-53 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5248 N$10496 N$10495 "Straight Waveguide" sch_x=-53 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5249 N$10498 N$10497 "Straight Waveguide" sch_x=-53 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5250 N$10500 N$10499 "Straight Waveguide" sch_x=-53 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5251 N$10502 N$10501 "Straight Waveguide" sch_x=-51 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5252 N$10504 N$10503 "Straight Waveguide" sch_x=-51 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5253 N$10506 N$10505 "Straight Waveguide" sch_x=-51 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5254 N$10508 N$10507 "Straight Waveguide" sch_x=-51 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5255 N$10510 N$10509 "Straight Waveguide" sch_x=-51 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5256 N$10512 N$10511 "Straight Waveguide" sch_x=-51 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5257 N$10514 N$10513 "Straight Waveguide" sch_x=-51 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5258 N$10516 N$10515 "Straight Waveguide" sch_x=-51 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5259 N$10518 N$10517 "Straight Waveguide" sch_x=-51 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5260 N$10520 N$10519 "Straight Waveguide" sch_x=-51 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5261 N$10522 N$10521 "Straight Waveguide" sch_x=-51 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5262 N$10524 N$10523 "Straight Waveguide" sch_x=-51 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5263 N$10526 N$10525 "Straight Waveguide" sch_x=-51 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5264 N$10528 N$10527 "Straight Waveguide" sch_x=-51 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5265 N$10530 N$10529 "Straight Waveguide" sch_x=-51 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5266 N$10532 N$10531 "Straight Waveguide" sch_x=-51 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5267 N$10534 N$10533 "Straight Waveguide" sch_x=-51 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5268 N$10536 N$10535 "Straight Waveguide" sch_x=-51 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5269 N$10538 N$10537 "Straight Waveguide" sch_x=-51 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5270 N$10540 N$10539 "Straight Waveguide" sch_x=-51 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5271 N$10542 N$10541 "Straight Waveguide" sch_x=-49 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5272 N$10544 N$10543 "Straight Waveguide" sch_x=-49 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5273 N$10546 N$10545 "Straight Waveguide" sch_x=-49 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5274 N$10548 N$10547 "Straight Waveguide" sch_x=-49 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5275 N$10550 N$10549 "Straight Waveguide" sch_x=-49 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5276 N$10552 N$10551 "Straight Waveguide" sch_x=-49 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5277 N$10554 N$10553 "Straight Waveguide" sch_x=-49 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5278 N$10556 N$10555 "Straight Waveguide" sch_x=-49 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5279 N$10558 N$10557 "Straight Waveguide" sch_x=-49 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5280 N$10560 N$10559 "Straight Waveguide" sch_x=-49 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5281 N$10562 N$10561 "Straight Waveguide" sch_x=-49 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5282 N$10564 N$10563 "Straight Waveguide" sch_x=-49 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5283 N$10566 N$10565 "Straight Waveguide" sch_x=-49 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5284 N$10568 N$10567 "Straight Waveguide" sch_x=-49 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5285 N$10570 N$10569 "Straight Waveguide" sch_x=-49 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5286 N$10572 N$10571 "Straight Waveguide" sch_x=-49 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5287 N$10574 N$10573 "Straight Waveguide" sch_x=-49 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5288 N$10576 N$10575 "Straight Waveguide" sch_x=-49 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5289 N$10578 N$10577 "Straight Waveguide" sch_x=-47 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5290 N$10580 N$10579 "Straight Waveguide" sch_x=-47 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5291 N$10582 N$10581 "Straight Waveguide" sch_x=-47 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5292 N$10584 N$10583 "Straight Waveguide" sch_x=-47 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5293 N$10586 N$10585 "Straight Waveguide" sch_x=-47 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5294 N$10588 N$10587 "Straight Waveguide" sch_x=-47 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5295 N$10590 N$10589 "Straight Waveguide" sch_x=-47 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5296 N$10592 N$10591 "Straight Waveguide" sch_x=-47 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5297 N$10594 N$10593 "Straight Waveguide" sch_x=-47 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5298 N$10596 N$10595 "Straight Waveguide" sch_x=-47 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5299 N$10598 N$10597 "Straight Waveguide" sch_x=-47 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5300 N$10600 N$10599 "Straight Waveguide" sch_x=-47 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5301 N$10602 N$10601 "Straight Waveguide" sch_x=-47 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5302 N$10604 N$10603 "Straight Waveguide" sch_x=-47 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5303 N$10606 N$10605 "Straight Waveguide" sch_x=-47 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5304 N$10608 N$10607 "Straight Waveguide" sch_x=-47 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5305 N$10610 N$10609 "Straight Waveguide" sch_x=-45 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5306 N$10612 N$10611 "Straight Waveguide" sch_x=-45 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5307 N$10614 N$10613 "Straight Waveguide" sch_x=-45 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5308 N$10616 N$10615 "Straight Waveguide" sch_x=-45 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5309 N$10618 N$10617 "Straight Waveguide" sch_x=-45 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5310 N$10620 N$10619 "Straight Waveguide" sch_x=-45 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5311 N$10622 N$10621 "Straight Waveguide" sch_x=-45 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5312 N$10624 N$10623 "Straight Waveguide" sch_x=-45 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5313 N$10626 N$10625 "Straight Waveguide" sch_x=-45 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5314 N$10628 N$10627 "Straight Waveguide" sch_x=-45 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5315 N$10630 N$10629 "Straight Waveguide" sch_x=-45 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5316 N$10632 N$10631 "Straight Waveguide" sch_x=-45 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5317 N$10634 N$10633 "Straight Waveguide" sch_x=-45 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5318 N$10636 N$10635 "Straight Waveguide" sch_x=-45 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5319 N$10638 N$10637 "Straight Waveguide" sch_x=-43 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5320 N$10640 N$10639 "Straight Waveguide" sch_x=-43 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5321 N$10642 N$10641 "Straight Waveguide" sch_x=-43 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5322 N$10644 N$10643 "Straight Waveguide" sch_x=-43 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5323 N$10646 N$10645 "Straight Waveguide" sch_x=-43 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5324 N$10648 N$10647 "Straight Waveguide" sch_x=-43 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5325 N$10650 N$10649 "Straight Waveguide" sch_x=-43 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5326 N$10652 N$10651 "Straight Waveguide" sch_x=-43 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5327 N$10654 N$10653 "Straight Waveguide" sch_x=-43 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5328 N$10656 N$10655 "Straight Waveguide" sch_x=-43 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5329 N$10658 N$10657 "Straight Waveguide" sch_x=-43 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5330 N$10660 N$10659 "Straight Waveguide" sch_x=-43 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5331 N$10662 N$10661 "Straight Waveguide" sch_x=-41 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5332 N$10664 N$10663 "Straight Waveguide" sch_x=-41 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5333 N$10666 N$10665 "Straight Waveguide" sch_x=-41 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5334 N$10668 N$10667 "Straight Waveguide" sch_x=-41 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5335 N$10670 N$10669 "Straight Waveguide" sch_x=-41 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5336 N$10672 N$10671 "Straight Waveguide" sch_x=-41 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5337 N$10674 N$10673 "Straight Waveguide" sch_x=-41 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5338 N$10676 N$10675 "Straight Waveguide" sch_x=-41 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5339 N$10678 N$10677 "Straight Waveguide" sch_x=-41 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5340 N$10680 N$10679 "Straight Waveguide" sch_x=-41 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5341 N$10682 N$10681 "Straight Waveguide" sch_x=-39 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5342 N$10684 N$10683 "Straight Waveguide" sch_x=-39 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5343 N$10686 N$10685 "Straight Waveguide" sch_x=-39 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5344 N$10688 N$10687 "Straight Waveguide" sch_x=-39 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5345 N$10690 N$10689 "Straight Waveguide" sch_x=-39 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5346 N$10692 N$10691 "Straight Waveguide" sch_x=-39 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5347 N$10694 N$10693 "Straight Waveguide" sch_x=-39 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5348 N$10696 N$10695 "Straight Waveguide" sch_x=-39 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5349 N$10698 N$10697 "Straight Waveguide" sch_x=-37 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5350 N$10700 N$10699 "Straight Waveguide" sch_x=-37 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5351 N$10702 N$10701 "Straight Waveguide" sch_x=-37 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5352 N$10704 N$10703 "Straight Waveguide" sch_x=-37 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5353 N$10706 N$10705 "Straight Waveguide" sch_x=-37 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5354 N$10708 N$10707 "Straight Waveguide" sch_x=-37 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5355 N$10710 N$10709 "Straight Waveguide" sch_x=-35 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5356 N$10712 N$10711 "Straight Waveguide" sch_x=-35 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5357 N$10714 N$10713 "Straight Waveguide" sch_x=-35 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5358 N$10716 N$10715 "Straight Waveguide" sch_x=-35 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5359 N$10718 N$10717 "Straight Waveguide" sch_x=-33 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5360 N$10720 N$10719 "Straight Waveguide" sch_x=-33 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5361 N$10721 N$10722 "Straight Waveguide" sch_x=-45 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5362 N$10723 N$10724 "Straight Waveguide" sch_x=-44 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5363 N$10725 N$10726 "Straight Waveguide" sch_x=-43 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5364 N$10727 N$10728 "Straight Waveguide" sch_x=-42 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5365 N$10729 N$10730 "Straight Waveguide" sch_x=-41 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5366 N$10731 N$10732 "Straight Waveguide" sch_x=-40 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5367 N$10733 N$10734 "Straight Waveguide" sch_x=-39 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5368 N$10735 N$10736 "Straight Waveguide" sch_x=-38 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5369 N$10737 N$10738 "Straight Waveguide" sch_x=-37 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5370 N$10739 N$10740 "Straight Waveguide" sch_x=-36 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5371 N$10741 N$10742 "Straight Waveguide" sch_x=-35 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5372 N$10743 N$10744 "Straight Waveguide" sch_x=-34 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5373 N$10745 N$10746 "Straight Waveguide" sch_x=-33 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5374 N$10747 N$10748 "Straight Waveguide" sch_x=-32 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5375 N$10749 N$10750 "Straight Waveguide" sch_x=-31 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5376 N$10751 N$10752 "Straight Waveguide" sch_x=-31 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5377 N$10753 N$10754 "Straight Waveguide" sch_x=-32 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5378 N$10755 N$10756 "Straight Waveguide" sch_x=-33 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5379 N$10757 N$10758 "Straight Waveguide" sch_x=-34 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5380 N$10759 N$10760 "Straight Waveguide" sch_x=-35 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5381 N$10761 N$10762 "Straight Waveguide" sch_x=-36 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5382 N$10763 N$10764 "Straight Waveguide" sch_x=-37 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5383 N$10765 N$10766 "Straight Waveguide" sch_x=-38 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5384 N$10767 N$10768 "Straight Waveguide" sch_x=-39 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5385 N$10769 N$10770 "Straight Waveguide" sch_x=-40 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5386 N$10771 N$10772 "Straight Waveguide" sch_x=-41 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5387 N$10773 N$10774 "Straight Waveguide" sch_x=-42 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5388 N$10775 N$10776 "Straight Waveguide" sch_x=-43 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5389 N$10777 N$10778 "Straight Waveguide" sch_x=-44 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5390 N$10779 N$10780 "Straight Waveguide" sch_x=-45 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5391 N$10781 N$10782 "Straight Waveguide" sch_x=-46 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5392 N$10783 N$10784 "Straight Waveguide" sch_x=-46 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5393 N$10785 N$10786 "Straight Waveguide" sch_x=61 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5394 N$10787 N$10788 "Straight Waveguide" sch_x=61 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5395 N$10789 N$10790 "Straight Waveguide" sch_x=61 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5396 N$10791 N$10792 "Straight Waveguide" sch_x=61 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5397 N$10793 N$10794 "Straight Waveguide" sch_x=61 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5398 N$10795 N$10796 "Straight Waveguide" sch_x=61 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5399 N$10797 N$10798 "Straight Waveguide" sch_x=61 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5400 N$10799 N$10800 "Straight Waveguide" sch_x=61 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5401 N$10801 N$10802 "Straight Waveguide" sch_x=61 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5402 N$10803 N$10804 "Straight Waveguide" sch_x=61 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5403 N$10805 N$10806 "Straight Waveguide" sch_x=61 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5404 N$10807 N$10808 "Straight Waveguide" sch_x=61 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5405 N$10809 N$10810 "Straight Waveguide" sch_x=61 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5406 N$10811 N$10812 "Straight Waveguide" sch_x=61 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5407 N$10813 N$10814 "Straight Waveguide" sch_x=61 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5408 N$10815 N$10816 "Straight Waveguide" sch_x=61 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5409 N$10817 N$10818 "Straight Waveguide" sch_x=61 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5410 N$10819 N$10820 "Straight Waveguide" sch_x=61 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5411 N$10821 N$10822 "Straight Waveguide" sch_x=61 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5412 N$10823 N$10824 "Straight Waveguide" sch_x=61 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5413 N$10825 N$10826 "Straight Waveguide" sch_x=61 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5414 N$10827 N$10828 "Straight Waveguide" sch_x=61 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5415 N$10829 N$10830 "Straight Waveguide" sch_x=61 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5416 N$10831 N$10832 "Straight Waveguide" sch_x=61 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5417 N$10833 N$10834 "Straight Waveguide" sch_x=61 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5418 N$10835 N$10836 "Straight Waveguide" sch_x=61 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5419 N$10837 N$10838 "Straight Waveguide" sch_x=61 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5420 N$10839 N$10840 "Straight Waveguide" sch_x=61 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5421 N$10841 N$10842 "Straight Waveguide" sch_x=61 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5422 N$10843 N$10844 "Straight Waveguide" sch_x=61 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5423 N$10845 N$10846 "Straight Waveguide" sch_x=59 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5424 N$10847 N$10848 "Straight Waveguide" sch_x=59 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5425 N$10849 N$10850 "Straight Waveguide" sch_x=59 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5426 N$10851 N$10852 "Straight Waveguide" sch_x=59 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5427 N$10853 N$10854 "Straight Waveguide" sch_x=59 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5428 N$10855 N$10856 "Straight Waveguide" sch_x=59 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5429 N$10857 N$10858 "Straight Waveguide" sch_x=59 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5430 N$10859 N$10860 "Straight Waveguide" sch_x=59 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5431 N$10861 N$10862 "Straight Waveguide" sch_x=59 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5432 N$10863 N$10864 "Straight Waveguide" sch_x=59 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5433 N$10865 N$10866 "Straight Waveguide" sch_x=59 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5434 N$10867 N$10868 "Straight Waveguide" sch_x=59 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5435 N$10869 N$10870 "Straight Waveguide" sch_x=59 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5436 N$10871 N$10872 "Straight Waveguide" sch_x=59 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5437 N$10873 N$10874 "Straight Waveguide" sch_x=59 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5438 N$10875 N$10876 "Straight Waveguide" sch_x=59 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5439 N$10877 N$10878 "Straight Waveguide" sch_x=59 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5440 N$10879 N$10880 "Straight Waveguide" sch_x=59 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5441 N$10881 N$10882 "Straight Waveguide" sch_x=59 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5442 N$10883 N$10884 "Straight Waveguide" sch_x=59 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5443 N$10885 N$10886 "Straight Waveguide" sch_x=59 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5444 N$10887 N$10888 "Straight Waveguide" sch_x=59 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5445 N$10889 N$10890 "Straight Waveguide" sch_x=59 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5446 N$10891 N$10892 "Straight Waveguide" sch_x=59 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5447 N$10893 N$10894 "Straight Waveguide" sch_x=59 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5448 N$10895 N$10896 "Straight Waveguide" sch_x=59 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5449 N$10897 N$10898 "Straight Waveguide" sch_x=59 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5450 N$10899 N$10900 "Straight Waveguide" sch_x=59 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5451 N$10901 N$10902 "Straight Waveguide" sch_x=57 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5452 N$10903 N$10904 "Straight Waveguide" sch_x=57 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5453 N$10905 N$10906 "Straight Waveguide" sch_x=57 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5454 N$10907 N$10908 "Straight Waveguide" sch_x=57 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5455 N$10909 N$10910 "Straight Waveguide" sch_x=57 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5456 N$10911 N$10912 "Straight Waveguide" sch_x=57 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5457 N$10913 N$10914 "Straight Waveguide" sch_x=57 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5458 N$10915 N$10916 "Straight Waveguide" sch_x=57 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5459 N$10917 N$10918 "Straight Waveguide" sch_x=57 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5460 N$10919 N$10920 "Straight Waveguide" sch_x=57 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5461 N$10921 N$10922 "Straight Waveguide" sch_x=57 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5462 N$10923 N$10924 "Straight Waveguide" sch_x=57 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5463 N$10925 N$10926 "Straight Waveguide" sch_x=57 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5464 N$10927 N$10928 "Straight Waveguide" sch_x=57 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5465 N$10929 N$10930 "Straight Waveguide" sch_x=57 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5466 N$10931 N$10932 "Straight Waveguide" sch_x=57 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5467 N$10933 N$10934 "Straight Waveguide" sch_x=57 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5468 N$10935 N$10936 "Straight Waveguide" sch_x=57 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5469 N$10937 N$10938 "Straight Waveguide" sch_x=57 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5470 N$10939 N$10940 "Straight Waveguide" sch_x=57 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5471 N$10941 N$10942 "Straight Waveguide" sch_x=57 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5472 N$10943 N$10944 "Straight Waveguide" sch_x=57 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5473 N$10945 N$10946 "Straight Waveguide" sch_x=57 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5474 N$10947 N$10948 "Straight Waveguide" sch_x=57 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5475 N$10949 N$10950 "Straight Waveguide" sch_x=57 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5476 N$10951 N$10952 "Straight Waveguide" sch_x=57 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5477 N$10953 N$10954 "Straight Waveguide" sch_x=55 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5478 N$10955 N$10956 "Straight Waveguide" sch_x=55 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5479 N$10957 N$10958 "Straight Waveguide" sch_x=55 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5480 N$10959 N$10960 "Straight Waveguide" sch_x=55 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5481 N$10961 N$10962 "Straight Waveguide" sch_x=55 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5482 N$10963 N$10964 "Straight Waveguide" sch_x=55 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5483 N$10965 N$10966 "Straight Waveguide" sch_x=55 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5484 N$10967 N$10968 "Straight Waveguide" sch_x=55 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5485 N$10969 N$10970 "Straight Waveguide" sch_x=55 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5486 N$10971 N$10972 "Straight Waveguide" sch_x=55 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5487 N$10973 N$10974 "Straight Waveguide" sch_x=55 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5488 N$10975 N$10976 "Straight Waveguide" sch_x=55 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5489 N$10977 N$10978 "Straight Waveguide" sch_x=55 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5490 N$10979 N$10980 "Straight Waveguide" sch_x=55 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5491 N$10981 N$10982 "Straight Waveguide" sch_x=55 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5492 N$10983 N$10984 "Straight Waveguide" sch_x=55 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5493 N$10985 N$10986 "Straight Waveguide" sch_x=55 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5494 N$10987 N$10988 "Straight Waveguide" sch_x=55 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5495 N$10989 N$10990 "Straight Waveguide" sch_x=55 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5496 N$10991 N$10992 "Straight Waveguide" sch_x=55 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5497 N$10993 N$10994 "Straight Waveguide" sch_x=55 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5498 N$10995 N$10996 "Straight Waveguide" sch_x=55 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5499 N$10997 N$10998 "Straight Waveguide" sch_x=55 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5500 N$10999 N$11000 "Straight Waveguide" sch_x=55 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5501 N$11001 N$11002 "Straight Waveguide" sch_x=53 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5502 N$11003 N$11004 "Straight Waveguide" sch_x=53 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5503 N$11005 N$11006 "Straight Waveguide" sch_x=53 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5504 N$11007 N$11008 "Straight Waveguide" sch_x=53 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5505 N$11009 N$11010 "Straight Waveguide" sch_x=53 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5506 N$11011 N$11012 "Straight Waveguide" sch_x=53 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5507 N$11013 N$11014 "Straight Waveguide" sch_x=53 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5508 N$11015 N$11016 "Straight Waveguide" sch_x=53 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5509 N$11017 N$11018 "Straight Waveguide" sch_x=53 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5510 N$11019 N$11020 "Straight Waveguide" sch_x=53 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5511 N$11021 N$11022 "Straight Waveguide" sch_x=53 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5512 N$11023 N$11024 "Straight Waveguide" sch_x=53 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5513 N$11025 N$11026 "Straight Waveguide" sch_x=53 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5514 N$11027 N$11028 "Straight Waveguide" sch_x=53 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5515 N$11029 N$11030 "Straight Waveguide" sch_x=53 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5516 N$11031 N$11032 "Straight Waveguide" sch_x=53 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5517 N$11033 N$11034 "Straight Waveguide" sch_x=53 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5518 N$11035 N$11036 "Straight Waveguide" sch_x=53 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5519 N$11037 N$11038 "Straight Waveguide" sch_x=53 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5520 N$11039 N$11040 "Straight Waveguide" sch_x=53 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5521 N$11041 N$11042 "Straight Waveguide" sch_x=53 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5522 N$11043 N$11044 "Straight Waveguide" sch_x=53 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5523 N$11045 N$11046 "Straight Waveguide" sch_x=51 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5524 N$11047 N$11048 "Straight Waveguide" sch_x=51 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5525 N$11049 N$11050 "Straight Waveguide" sch_x=51 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5526 N$11051 N$11052 "Straight Waveguide" sch_x=51 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5527 N$11053 N$11054 "Straight Waveguide" sch_x=51 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5528 N$11055 N$11056 "Straight Waveguide" sch_x=51 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5529 N$11057 N$11058 "Straight Waveguide" sch_x=51 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5530 N$11059 N$11060 "Straight Waveguide" sch_x=51 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5531 N$11061 N$11062 "Straight Waveguide" sch_x=51 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5532 N$11063 N$11064 "Straight Waveguide" sch_x=51 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5533 N$11065 N$11066 "Straight Waveguide" sch_x=51 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5534 N$11067 N$11068 "Straight Waveguide" sch_x=51 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5535 N$11069 N$11070 "Straight Waveguide" sch_x=51 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5536 N$11071 N$11072 "Straight Waveguide" sch_x=51 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5537 N$11073 N$11074 "Straight Waveguide" sch_x=51 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5538 N$11075 N$11076 "Straight Waveguide" sch_x=51 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5539 N$11077 N$11078 "Straight Waveguide" sch_x=51 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5540 N$11079 N$11080 "Straight Waveguide" sch_x=51 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5541 N$11081 N$11082 "Straight Waveguide" sch_x=51 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5542 N$11083 N$11084 "Straight Waveguide" sch_x=51 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5543 N$11085 N$11086 "Straight Waveguide" sch_x=49 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5544 N$11087 N$11088 "Straight Waveguide" sch_x=49 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5545 N$11089 N$11090 "Straight Waveguide" sch_x=49 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5546 N$11091 N$11092 "Straight Waveguide" sch_x=49 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5547 N$11093 N$11094 "Straight Waveguide" sch_x=49 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5548 N$11095 N$11096 "Straight Waveguide" sch_x=49 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5549 N$11097 N$11098 "Straight Waveguide" sch_x=49 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5550 N$11099 N$11100 "Straight Waveguide" sch_x=49 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5551 N$11101 N$11102 "Straight Waveguide" sch_x=49 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5552 N$11103 N$11104 "Straight Waveguide" sch_x=49 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5553 N$11105 N$11106 "Straight Waveguide" sch_x=49 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5554 N$11107 N$11108 "Straight Waveguide" sch_x=49 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5555 N$11109 N$11110 "Straight Waveguide" sch_x=49 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5556 N$11111 N$11112 "Straight Waveguide" sch_x=49 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5557 N$11113 N$11114 "Straight Waveguide" sch_x=49 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5558 N$11115 N$11116 "Straight Waveguide" sch_x=49 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5559 N$11117 N$11118 "Straight Waveguide" sch_x=49 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5560 N$11119 N$11120 "Straight Waveguide" sch_x=49 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5561 N$11121 N$11122 "Straight Waveguide" sch_x=47 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5562 N$11123 N$11124 "Straight Waveguide" sch_x=47 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5563 N$11125 N$11126 "Straight Waveguide" sch_x=47 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5564 N$11127 N$11128 "Straight Waveguide" sch_x=47 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5565 N$11129 N$11130 "Straight Waveguide" sch_x=47 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5566 N$11131 N$11132 "Straight Waveguide" sch_x=47 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5567 N$11133 N$11134 "Straight Waveguide" sch_x=47 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5568 N$11135 N$11136 "Straight Waveguide" sch_x=47 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5569 N$11137 N$11138 "Straight Waveguide" sch_x=47 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5570 N$11139 N$11140 "Straight Waveguide" sch_x=47 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5571 N$11141 N$11142 "Straight Waveguide" sch_x=47 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5572 N$11143 N$11144 "Straight Waveguide" sch_x=47 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5573 N$11145 N$11146 "Straight Waveguide" sch_x=47 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5574 N$11147 N$11148 "Straight Waveguide" sch_x=47 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5575 N$11149 N$11150 "Straight Waveguide" sch_x=47 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5576 N$11151 N$11152 "Straight Waveguide" sch_x=47 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5577 N$11153 N$11154 "Straight Waveguide" sch_x=45 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5578 N$11155 N$11156 "Straight Waveguide" sch_x=45 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5579 N$11157 N$11158 "Straight Waveguide" sch_x=45 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5580 N$11159 N$11160 "Straight Waveguide" sch_x=45 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5581 N$11161 N$11162 "Straight Waveguide" sch_x=45 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5582 N$11163 N$11164 "Straight Waveguide" sch_x=45 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5583 N$11165 N$11166 "Straight Waveguide" sch_x=45 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5584 N$11167 N$11168 "Straight Waveguide" sch_x=45 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5585 N$11169 N$11170 "Straight Waveguide" sch_x=45 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5586 N$11171 N$11172 "Straight Waveguide" sch_x=45 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5587 N$11173 N$11174 "Straight Waveguide" sch_x=45 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5588 N$11175 N$11176 "Straight Waveguide" sch_x=45 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5589 N$11177 N$11178 "Straight Waveguide" sch_x=45 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5590 N$11179 N$11180 "Straight Waveguide" sch_x=45 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5591 N$11181 N$11182 "Straight Waveguide" sch_x=43 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5592 N$11183 N$11184 "Straight Waveguide" sch_x=43 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5593 N$11185 N$11186 "Straight Waveguide" sch_x=43 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5594 N$11187 N$11188 "Straight Waveguide" sch_x=43 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5595 N$11189 N$11190 "Straight Waveguide" sch_x=43 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5596 N$11191 N$11192 "Straight Waveguide" sch_x=43 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5597 N$11193 N$11194 "Straight Waveguide" sch_x=43 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5598 N$11195 N$11196 "Straight Waveguide" sch_x=43 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5599 N$11197 N$11198 "Straight Waveguide" sch_x=43 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5600 N$11199 N$11200 "Straight Waveguide" sch_x=43 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5601 N$11201 N$11202 "Straight Waveguide" sch_x=43 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5602 N$11203 N$11204 "Straight Waveguide" sch_x=43 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5603 N$11205 N$11206 "Straight Waveguide" sch_x=41 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5604 N$11207 N$11208 "Straight Waveguide" sch_x=41 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5605 N$11209 N$11210 "Straight Waveguide" sch_x=41 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5606 N$11211 N$11212 "Straight Waveguide" sch_x=41 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5607 N$11213 N$11214 "Straight Waveguide" sch_x=41 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5608 N$11215 N$11216 "Straight Waveguide" sch_x=41 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5609 N$11217 N$11218 "Straight Waveguide" sch_x=41 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5610 N$11219 N$11220 "Straight Waveguide" sch_x=41 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5611 N$11221 N$11222 "Straight Waveguide" sch_x=41 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5612 N$11223 N$11224 "Straight Waveguide" sch_x=41 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5613 N$11225 N$11226 "Straight Waveguide" sch_x=39 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5614 N$11227 N$11228 "Straight Waveguide" sch_x=39 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5615 N$11229 N$11230 "Straight Waveguide" sch_x=39 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5616 N$11231 N$11232 "Straight Waveguide" sch_x=39 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5617 N$11233 N$11234 "Straight Waveguide" sch_x=39 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5618 N$11235 N$11236 "Straight Waveguide" sch_x=39 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5619 N$11237 N$11238 "Straight Waveguide" sch_x=39 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5620 N$11239 N$11240 "Straight Waveguide" sch_x=39 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5621 N$11241 N$11242 "Straight Waveguide" sch_x=37 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5622 N$11243 N$11244 "Straight Waveguide" sch_x=37 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5623 N$11245 N$11246 "Straight Waveguide" sch_x=37 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5624 N$11247 N$11248 "Straight Waveguide" sch_x=37 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5625 N$11249 N$11250 "Straight Waveguide" sch_x=37 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5626 N$11251 N$11252 "Straight Waveguide" sch_x=37 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5627 N$11253 N$11254 "Straight Waveguide" sch_x=35 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5628 N$11255 N$11256 "Straight Waveguide" sch_x=35 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5629 N$11257 N$11258 "Straight Waveguide" sch_x=35 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5630 N$11259 N$11260 "Straight Waveguide" sch_x=35 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5631 N$11261 N$11262 "Straight Waveguide" sch_x=33 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5632 N$11263 N$11264 "Straight Waveguide" sch_x=33 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5633 N$11266 N$11265 "Straight Waveguide" sch_x=45 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5634 N$11268 N$11267 "Straight Waveguide" sch_x=44 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5635 N$11270 N$11269 "Straight Waveguide" sch_x=43 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5636 N$11272 N$11271 "Straight Waveguide" sch_x=42 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5637 N$11274 N$11273 "Straight Waveguide" sch_x=41 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5638 N$11276 N$11275 "Straight Waveguide" sch_x=40 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5639 N$11278 N$11277 "Straight Waveguide" sch_x=39 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5640 N$11280 N$11279 "Straight Waveguide" sch_x=38 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5641 N$11282 N$11281 "Straight Waveguide" sch_x=37 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5642 N$11284 N$11283 "Straight Waveguide" sch_x=36 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5643 N$11286 N$11285 "Straight Waveguide" sch_x=35 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5644 N$11288 N$11287 "Straight Waveguide" sch_x=34 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5645 N$11290 N$11289 "Straight Waveguide" sch_x=33 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5646 N$11292 N$11291 "Straight Waveguide" sch_x=32 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5647 N$11294 N$11293 "Straight Waveguide" sch_x=31 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5648 N$11296 N$11295 "Straight Waveguide" sch_x=31 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5649 N$11298 N$11297 "Straight Waveguide" sch_x=32 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5650 N$11300 N$11299 "Straight Waveguide" sch_x=33 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5651 N$11302 N$11301 "Straight Waveguide" sch_x=34 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5652 N$11304 N$11303 "Straight Waveguide" sch_x=35 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5653 N$11306 N$11305 "Straight Waveguide" sch_x=36 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5654 N$11308 N$11307 "Straight Waveguide" sch_x=37 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5655 N$11310 N$11309 "Straight Waveguide" sch_x=38 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5656 N$11312 N$11311 "Straight Waveguide" sch_x=39 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5657 N$11314 N$11313 "Straight Waveguide" sch_x=40 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5658 N$11316 N$11315 "Straight Waveguide" sch_x=41 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5659 N$11318 N$11317 "Straight Waveguide" sch_x=42 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5660 N$11320 N$11319 "Straight Waveguide" sch_x=43 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5661 N$11322 N$11321 "Straight Waveguide" sch_x=44 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5662 N$11324 N$11323 "Straight Waveguide" sch_x=45 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5663 N$11326 N$11325 "Straight Waveguide" sch_x=46 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5664 N$11328 N$11327 "Straight Waveguide" sch_x=46 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5665 N$11329 N$11330 "Straight Waveguide" sch_x=-4 sch_y=-32.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5666 N$11331 N$11332 "Straight Waveguide" sch_x=-5 sch_y=-33.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5667 N$11333 N$11334 "Straight Waveguide" sch_x=-5 sch_y=-34.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5668 N$11335 N$11336 "Straight Waveguide" sch_x=-3 sch_y=-33.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5669 N$11337 N$11338 "Straight Waveguide" sch_x=-3 sch_y=-34.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5670 N$11339 N$11340 "Straight Waveguide" sch_x=-4 sch_y=-35.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5671 N$11341 N$11342 "Straight Waveguide" sch_x=0 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5672 N$11343 N$11344 "Straight Waveguide" sch_x=-1 sch_y=-32.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5673 N$11345 N$11346 "Straight Waveguide" sch_x=-1 sch_y=-33.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5674 N$11347 N$11348 "Straight Waveguide" sch_x=1 sch_y=-33.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5675 N$11349 N$11350 "Straight Waveguide" sch_x=1 sch_y=-32.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5676 N$11351 N$11352 "Straight Waveguide" sch_x=0 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5677 N$11353 N$11354 "Straight Waveguide" sch_x=0 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5678 N$11355 N$11356 "Straight Waveguide" sch_x=-1 sch_y=-34.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5679 N$11357 N$11358 "Straight Waveguide" sch_x=-1 sch_y=-35.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5680 N$11359 N$11360 "Straight Waveguide" sch_x=1 sch_y=-35.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5681 N$11361 N$11362 "Straight Waveguide" sch_x=1 sch_y=-34.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5682 N$11363 N$11364 "Straight Waveguide" sch_x=0 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5683 N$11365 N$11366 "Straight Waveguide" sch_x=4 sch_y=-32.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5684 N$11367 N$11368 "Straight Waveguide" sch_x=3 sch_y=-33.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5685 N$11369 N$11370 "Straight Waveguide" sch_x=3 sch_y=-34.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5686 N$11371 N$11372 "Straight Waveguide" sch_x=5 sch_y=-34.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5687 N$11373 N$11374 "Straight Waveguide" sch_x=5 sch_y=-33.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5688 N$11375 N$11376 "Straight Waveguide" sch_x=4 sch_y=-35.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5689 N$11377 N$11378 "Straight Waveguide" sch_x=-4 sch_y=-36.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5690 N$11379 N$11380 "Straight Waveguide" sch_x=-5 sch_y=-37.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5691 N$11381 N$11382 "Straight Waveguide" sch_x=-5 sch_y=-38.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5692 N$11383 N$11384 "Straight Waveguide" sch_x=-3 sch_y=-37.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5693 N$11385 N$11386 "Straight Waveguide" sch_x=-3 sch_y=-38.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5694 N$11387 N$11388 "Straight Waveguide" sch_x=-4 sch_y=-39.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5695 N$11389 N$11390 "Straight Waveguide" sch_x=0 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5696 N$11391 N$11392 "Straight Waveguide" sch_x=-1 sch_y=-36.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5697 N$11393 N$11394 "Straight Waveguide" sch_x=-1 sch_y=-37.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5698 N$11395 N$11396 "Straight Waveguide" sch_x=1 sch_y=-37.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5699 N$11397 N$11398 "Straight Waveguide" sch_x=1 sch_y=-36.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5700 N$11399 N$11400 "Straight Waveguide" sch_x=0 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5701 N$11401 N$11402 "Straight Waveguide" sch_x=0 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5702 N$11403 N$11404 "Straight Waveguide" sch_x=-1 sch_y=-38.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5703 N$11405 N$11406 "Straight Waveguide" sch_x=-1 sch_y=-39.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5704 N$11407 N$11408 "Straight Waveguide" sch_x=1 sch_y=-39.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5705 N$11409 N$11410 "Straight Waveguide" sch_x=1 sch_y=-38.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5706 N$11411 N$11412 "Straight Waveguide" sch_x=0 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5707 N$11413 N$11414 "Straight Waveguide" sch_x=4 sch_y=-36.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5708 N$11415 N$11416 "Straight Waveguide" sch_x=3 sch_y=-37.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5709 N$11417 N$11418 "Straight Waveguide" sch_x=3 sch_y=-38.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5710 N$11419 N$11420 "Straight Waveguide" sch_x=5 sch_y=-38.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5711 N$11421 N$11422 "Straight Waveguide" sch_x=5 sch_y=-37.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5712 N$11423 N$11424 "Straight Waveguide" sch_x=4 sch_y=-39.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5713 N$11426 N$11425 "Straight Waveguide" sch_x=-13 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5714 N$11428 N$11427 "Straight Waveguide" sch_x=-13 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5715 N$11430 N$11429 "Straight Waveguide" sch_x=-13 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5716 N$11432 N$11431 "Straight Waveguide" sch_x=-13 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5717 N$11434 N$11433 "Straight Waveguide" sch_x=-13 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5718 N$11436 N$11435 "Straight Waveguide" sch_x=-13 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5719 N$11438 N$11437 "Straight Waveguide" sch_x=-11 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5720 N$11440 N$11439 "Straight Waveguide" sch_x=-11 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5721 N$11442 N$11441 "Straight Waveguide" sch_x=-11 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5722 N$11444 N$11443 "Straight Waveguide" sch_x=-11 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5723 N$11446 N$11445 "Straight Waveguide" sch_x=-9 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5724 N$11448 N$11447 "Straight Waveguide" sch_x=-9 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5725 N$11449 N$11450 "Straight Waveguide" sch_x=-9 sch_y=-33.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5726 N$11451 N$11452 "Straight Waveguide" sch_x=-8 sch_y=-34.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5727 N$11453 N$11454 "Straight Waveguide" sch_x=-7 sch_y=-35.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5728 N$11455 N$11456 "Straight Waveguide" sch_x=-7 sch_y=-36.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5729 N$11457 N$11458 "Straight Waveguide" sch_x=-8 sch_y=-37.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5730 N$11459 N$11460 "Straight Waveguide" sch_x=-9 sch_y=-38.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5731 N$11461 N$11462 "Straight Waveguide" sch_x=-10 sch_y=-33.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5732 N$11463 N$11464 "Straight Waveguide" sch_x=-10 sch_y=-38.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5733 N$11465 N$11466 "Straight Waveguide" sch_x=13 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5734 N$11467 N$11468 "Straight Waveguide" sch_x=13 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5735 N$11469 N$11470 "Straight Waveguide" sch_x=13 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5736 N$11471 N$11472 "Straight Waveguide" sch_x=13 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5737 N$11473 N$11474 "Straight Waveguide" sch_x=13 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5738 N$11475 N$11476 "Straight Waveguide" sch_x=13 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5739 N$11477 N$11478 "Straight Waveguide" sch_x=11 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5740 N$11479 N$11480 "Straight Waveguide" sch_x=11 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5741 N$11481 N$11482 "Straight Waveguide" sch_x=11 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5742 N$11483 N$11484 "Straight Waveguide" sch_x=11 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5743 N$11485 N$11486 "Straight Waveguide" sch_x=9 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5744 N$11487 N$11488 "Straight Waveguide" sch_x=9 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5745 N$11490 N$11489 "Straight Waveguide" sch_x=9 sch_y=-33.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5746 N$11492 N$11491 "Straight Waveguide" sch_x=8 sch_y=-34.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5747 N$11494 N$11493 "Straight Waveguide" sch_x=7 sch_y=-35.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5748 N$11496 N$11495 "Straight Waveguide" sch_x=7 sch_y=-36.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5749 N$11498 N$11497 "Straight Waveguide" sch_x=8 sch_y=-37.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5750 N$11500 N$11499 "Straight Waveguide" sch_x=9 sch_y=-38.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5751 N$11502 N$11501 "Straight Waveguide" sch_x=10 sch_y=-33.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5752 N$11504 N$11503 "Straight Waveguide" sch_x=10 sch_y=-38.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5753 N$11505 N$11506 "Straight Waveguide" sch_x=-4 sch_y=-40.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5754 N$11507 N$11508 "Straight Waveguide" sch_x=-5 sch_y=-41.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5755 N$11509 N$11510 "Straight Waveguide" sch_x=-5 sch_y=-42.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5756 N$11511 N$11512 "Straight Waveguide" sch_x=-3 sch_y=-41.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5757 N$11513 N$11514 "Straight Waveguide" sch_x=-3 sch_y=-42.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5758 N$11515 N$11516 "Straight Waveguide" sch_x=-4 sch_y=-43.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5759 N$11517 N$11518 "Straight Waveguide" sch_x=0 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5760 N$11519 N$11520 "Straight Waveguide" sch_x=-1 sch_y=-40.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5761 N$11521 N$11522 "Straight Waveguide" sch_x=-1 sch_y=-41.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5762 N$11523 N$11524 "Straight Waveguide" sch_x=1 sch_y=-41.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5763 N$11525 N$11526 "Straight Waveguide" sch_x=1 sch_y=-40.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5764 N$11527 N$11528 "Straight Waveguide" sch_x=0 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5765 N$11529 N$11530 "Straight Waveguide" sch_x=0 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5766 N$11531 N$11532 "Straight Waveguide" sch_x=-1 sch_y=-42.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5767 N$11533 N$11534 "Straight Waveguide" sch_x=-1 sch_y=-43.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5768 N$11535 N$11536 "Straight Waveguide" sch_x=1 sch_y=-43.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5769 N$11537 N$11538 "Straight Waveguide" sch_x=1 sch_y=-42.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5770 N$11539 N$11540 "Straight Waveguide" sch_x=0 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5771 N$11541 N$11542 "Straight Waveguide" sch_x=4 sch_y=-40.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5772 N$11543 N$11544 "Straight Waveguide" sch_x=3 sch_y=-41.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5773 N$11545 N$11546 "Straight Waveguide" sch_x=3 sch_y=-42.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5774 N$11547 N$11548 "Straight Waveguide" sch_x=5 sch_y=-42.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5775 N$11549 N$11550 "Straight Waveguide" sch_x=5 sch_y=-41.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5776 N$11551 N$11552 "Straight Waveguide" sch_x=4 sch_y=-43.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5777 N$11553 N$11554 "Straight Waveguide" sch_x=-4 sch_y=-44.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5778 N$11555 N$11556 "Straight Waveguide" sch_x=-5 sch_y=-45.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5779 N$11557 N$11558 "Straight Waveguide" sch_x=-5 sch_y=-46.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5780 N$11559 N$11560 "Straight Waveguide" sch_x=-3 sch_y=-45.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5781 N$11561 N$11562 "Straight Waveguide" sch_x=-3 sch_y=-46.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5782 N$11563 N$11564 "Straight Waveguide" sch_x=-4 sch_y=-47.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5783 N$11565 N$11566 "Straight Waveguide" sch_x=0 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5784 N$11567 N$11568 "Straight Waveguide" sch_x=-1 sch_y=-44.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5785 N$11569 N$11570 "Straight Waveguide" sch_x=-1 sch_y=-45.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5786 N$11571 N$11572 "Straight Waveguide" sch_x=1 sch_y=-45.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5787 N$11573 N$11574 "Straight Waveguide" sch_x=1 sch_y=-44.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5788 N$11575 N$11576 "Straight Waveguide" sch_x=0 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5789 N$11577 N$11578 "Straight Waveguide" sch_x=0 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5790 N$11579 N$11580 "Straight Waveguide" sch_x=-1 sch_y=-46.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5791 N$11581 N$11582 "Straight Waveguide" sch_x=-1 sch_y=-47.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5792 N$11583 N$11584 "Straight Waveguide" sch_x=1 sch_y=-47.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5793 N$11585 N$11586 "Straight Waveguide" sch_x=1 sch_y=-46.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5794 N$11587 N$11588 "Straight Waveguide" sch_x=0 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5795 N$11589 N$11590 "Straight Waveguide" sch_x=4 sch_y=-44.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5796 N$11591 N$11592 "Straight Waveguide" sch_x=3 sch_y=-45.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5797 N$11593 N$11594 "Straight Waveguide" sch_x=3 sch_y=-46.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5798 N$11595 N$11596 "Straight Waveguide" sch_x=5 sch_y=-46.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5799 N$11597 N$11598 "Straight Waveguide" sch_x=5 sch_y=-45.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5800 N$11599 N$11600 "Straight Waveguide" sch_x=4 sch_y=-47.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5801 N$11602 N$11601 "Straight Waveguide" sch_x=-13 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5802 N$11604 N$11603 "Straight Waveguide" sch_x=-13 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5803 N$11606 N$11605 "Straight Waveguide" sch_x=-13 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5804 N$11608 N$11607 "Straight Waveguide" sch_x=-13 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5805 N$11610 N$11609 "Straight Waveguide" sch_x=-13 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5806 N$11612 N$11611 "Straight Waveguide" sch_x=-13 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5807 N$11614 N$11613 "Straight Waveguide" sch_x=-11 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5808 N$11616 N$11615 "Straight Waveguide" sch_x=-11 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5809 N$11618 N$11617 "Straight Waveguide" sch_x=-11 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5810 N$11620 N$11619 "Straight Waveguide" sch_x=-11 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5811 N$11622 N$11621 "Straight Waveguide" sch_x=-9 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5812 N$11624 N$11623 "Straight Waveguide" sch_x=-9 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5813 N$11625 N$11626 "Straight Waveguide" sch_x=-9 sch_y=-41.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5814 N$11627 N$11628 "Straight Waveguide" sch_x=-8 sch_y=-42.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5815 N$11629 N$11630 "Straight Waveguide" sch_x=-7 sch_y=-43.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5816 N$11631 N$11632 "Straight Waveguide" sch_x=-7 sch_y=-44.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5817 N$11633 N$11634 "Straight Waveguide" sch_x=-8 sch_y=-45.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5818 N$11635 N$11636 "Straight Waveguide" sch_x=-9 sch_y=-46.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5819 N$11637 N$11638 "Straight Waveguide" sch_x=-10 sch_y=-41.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5820 N$11639 N$11640 "Straight Waveguide" sch_x=-10 sch_y=-46.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5821 N$11641 N$11642 "Straight Waveguide" sch_x=13 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5822 N$11643 N$11644 "Straight Waveguide" sch_x=13 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5823 N$11645 N$11646 "Straight Waveguide" sch_x=13 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5824 N$11647 N$11648 "Straight Waveguide" sch_x=13 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5825 N$11649 N$11650 "Straight Waveguide" sch_x=13 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5826 N$11651 N$11652 "Straight Waveguide" sch_x=13 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5827 N$11653 N$11654 "Straight Waveguide" sch_x=11 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5828 N$11655 N$11656 "Straight Waveguide" sch_x=11 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5829 N$11657 N$11658 "Straight Waveguide" sch_x=11 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5830 N$11659 N$11660 "Straight Waveguide" sch_x=11 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5831 N$11661 N$11662 "Straight Waveguide" sch_x=9 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5832 N$11663 N$11664 "Straight Waveguide" sch_x=9 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5833 N$11666 N$11665 "Straight Waveguide" sch_x=9 sch_y=-41.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5834 N$11668 N$11667 "Straight Waveguide" sch_x=8 sch_y=-42.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5835 N$11670 N$11669 "Straight Waveguide" sch_x=7 sch_y=-43.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5836 N$11672 N$11671 "Straight Waveguide" sch_x=7 sch_y=-44.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5837 N$11674 N$11673 "Straight Waveguide" sch_x=8 sch_y=-45.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5838 N$11676 N$11675 "Straight Waveguide" sch_x=9 sch_y=-46.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5839 N$11678 N$11677 "Straight Waveguide" sch_x=10 sch_y=-41.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5840 N$11680 N$11679 "Straight Waveguide" sch_x=10 sch_y=-46.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5841 N$11682 N$11681 "Straight Waveguide" sch_x=-29 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5842 N$11684 N$11683 "Straight Waveguide" sch_x=-29 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5843 N$11686 N$11685 "Straight Waveguide" sch_x=-29 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5844 N$11688 N$11687 "Straight Waveguide" sch_x=-29 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5845 N$11690 N$11689 "Straight Waveguide" sch_x=-29 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5846 N$11692 N$11691 "Straight Waveguide" sch_x=-29 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5847 N$11694 N$11693 "Straight Waveguide" sch_x=-29 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5848 N$11696 N$11695 "Straight Waveguide" sch_x=-29 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5849 N$11698 N$11697 "Straight Waveguide" sch_x=-29 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5850 N$11700 N$11699 "Straight Waveguide" sch_x=-29 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5851 N$11702 N$11701 "Straight Waveguide" sch_x=-29 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5852 N$11704 N$11703 "Straight Waveguide" sch_x=-29 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5853 N$11706 N$11705 "Straight Waveguide" sch_x=-29 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5854 N$11708 N$11707 "Straight Waveguide" sch_x=-29 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5855 N$11710 N$11709 "Straight Waveguide" sch_x=-27 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5856 N$11712 N$11711 "Straight Waveguide" sch_x=-27 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5857 N$11714 N$11713 "Straight Waveguide" sch_x=-27 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5858 N$11716 N$11715 "Straight Waveguide" sch_x=-27 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5859 N$11718 N$11717 "Straight Waveguide" sch_x=-27 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5860 N$11720 N$11719 "Straight Waveguide" sch_x=-27 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5861 N$11722 N$11721 "Straight Waveguide" sch_x=-27 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5862 N$11724 N$11723 "Straight Waveguide" sch_x=-27 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5863 N$11726 N$11725 "Straight Waveguide" sch_x=-27 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5864 N$11728 N$11727 "Straight Waveguide" sch_x=-27 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5865 N$11730 N$11729 "Straight Waveguide" sch_x=-27 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5866 N$11732 N$11731 "Straight Waveguide" sch_x=-27 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5867 N$11734 N$11733 "Straight Waveguide" sch_x=-25 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5868 N$11736 N$11735 "Straight Waveguide" sch_x=-25 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5869 N$11738 N$11737 "Straight Waveguide" sch_x=-25 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5870 N$11740 N$11739 "Straight Waveguide" sch_x=-25 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5871 N$11742 N$11741 "Straight Waveguide" sch_x=-25 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5872 N$11744 N$11743 "Straight Waveguide" sch_x=-25 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5873 N$11746 N$11745 "Straight Waveguide" sch_x=-25 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5874 N$11748 N$11747 "Straight Waveguide" sch_x=-25 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5875 N$11750 N$11749 "Straight Waveguide" sch_x=-25 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5876 N$11752 N$11751 "Straight Waveguide" sch_x=-25 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5877 N$11754 N$11753 "Straight Waveguide" sch_x=-23 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5878 N$11756 N$11755 "Straight Waveguide" sch_x=-23 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5879 N$11758 N$11757 "Straight Waveguide" sch_x=-23 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5880 N$11760 N$11759 "Straight Waveguide" sch_x=-23 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5881 N$11762 N$11761 "Straight Waveguide" sch_x=-23 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5882 N$11764 N$11763 "Straight Waveguide" sch_x=-23 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5883 N$11766 N$11765 "Straight Waveguide" sch_x=-23 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5884 N$11768 N$11767 "Straight Waveguide" sch_x=-23 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5885 N$11770 N$11769 "Straight Waveguide" sch_x=-21 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5886 N$11772 N$11771 "Straight Waveguide" sch_x=-21 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5887 N$11774 N$11773 "Straight Waveguide" sch_x=-21 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5888 N$11776 N$11775 "Straight Waveguide" sch_x=-21 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5889 N$11778 N$11777 "Straight Waveguide" sch_x=-21 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5890 N$11780 N$11779 "Straight Waveguide" sch_x=-21 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5891 N$11782 N$11781 "Straight Waveguide" sch_x=-19 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5892 N$11784 N$11783 "Straight Waveguide" sch_x=-19 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5893 N$11786 N$11785 "Straight Waveguide" sch_x=-19 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5894 N$11788 N$11787 "Straight Waveguide" sch_x=-19 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5895 N$11790 N$11789 "Straight Waveguide" sch_x=-17 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5896 N$11792 N$11791 "Straight Waveguide" sch_x=-17 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5897 N$11793 N$11794 "Straight Waveguide" sch_x=-21 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5898 N$11795 N$11796 "Straight Waveguide" sch_x=-20 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5899 N$11797 N$11798 "Straight Waveguide" sch_x=-19 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5900 N$11799 N$11800 "Straight Waveguide" sch_x=-18 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5901 N$11801 N$11802 "Straight Waveguide" sch_x=-17 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5902 N$11803 N$11804 "Straight Waveguide" sch_x=-16 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5903 N$11805 N$11806 "Straight Waveguide" sch_x=-15 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5904 N$11807 N$11808 "Straight Waveguide" sch_x=-15 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5905 N$11809 N$11810 "Straight Waveguide" sch_x=-16 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5906 N$11811 N$11812 "Straight Waveguide" sch_x=-17 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5907 N$11813 N$11814 "Straight Waveguide" sch_x=-18 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5908 N$11815 N$11816 "Straight Waveguide" sch_x=-19 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5909 N$11817 N$11818 "Straight Waveguide" sch_x=-20 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5910 N$11819 N$11820 "Straight Waveguide" sch_x=-21 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5911 N$11821 N$11822 "Straight Waveguide" sch_x=-22 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5912 N$11823 N$11824 "Straight Waveguide" sch_x=-22 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5913 N$11825 N$11826 "Straight Waveguide" sch_x=29 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5914 N$11827 N$11828 "Straight Waveguide" sch_x=29 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5915 N$11829 N$11830 "Straight Waveguide" sch_x=29 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5916 N$11831 N$11832 "Straight Waveguide" sch_x=29 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5917 N$11833 N$11834 "Straight Waveguide" sch_x=29 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5918 N$11835 N$11836 "Straight Waveguide" sch_x=29 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5919 N$11837 N$11838 "Straight Waveguide" sch_x=29 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5920 N$11839 N$11840 "Straight Waveguide" sch_x=29 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5921 N$11841 N$11842 "Straight Waveguide" sch_x=29 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5922 N$11843 N$11844 "Straight Waveguide" sch_x=29 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5923 N$11845 N$11846 "Straight Waveguide" sch_x=29 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5924 N$11847 N$11848 "Straight Waveguide" sch_x=29 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5925 N$11849 N$11850 "Straight Waveguide" sch_x=29 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5926 N$11851 N$11852 "Straight Waveguide" sch_x=29 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5927 N$11853 N$11854 "Straight Waveguide" sch_x=27 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5928 N$11855 N$11856 "Straight Waveguide" sch_x=27 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5929 N$11857 N$11858 "Straight Waveguide" sch_x=27 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5930 N$11859 N$11860 "Straight Waveguide" sch_x=27 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5931 N$11861 N$11862 "Straight Waveguide" sch_x=27 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5932 N$11863 N$11864 "Straight Waveguide" sch_x=27 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5933 N$11865 N$11866 "Straight Waveguide" sch_x=27 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5934 N$11867 N$11868 "Straight Waveguide" sch_x=27 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5935 N$11869 N$11870 "Straight Waveguide" sch_x=27 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5936 N$11871 N$11872 "Straight Waveguide" sch_x=27 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5937 N$11873 N$11874 "Straight Waveguide" sch_x=27 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5938 N$11875 N$11876 "Straight Waveguide" sch_x=27 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5939 N$11877 N$11878 "Straight Waveguide" sch_x=25 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5940 N$11879 N$11880 "Straight Waveguide" sch_x=25 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5941 N$11881 N$11882 "Straight Waveguide" sch_x=25 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5942 N$11883 N$11884 "Straight Waveguide" sch_x=25 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5943 N$11885 N$11886 "Straight Waveguide" sch_x=25 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5944 N$11887 N$11888 "Straight Waveguide" sch_x=25 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5945 N$11889 N$11890 "Straight Waveguide" sch_x=25 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5946 N$11891 N$11892 "Straight Waveguide" sch_x=25 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5947 N$11893 N$11894 "Straight Waveguide" sch_x=25 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5948 N$11895 N$11896 "Straight Waveguide" sch_x=25 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5949 N$11897 N$11898 "Straight Waveguide" sch_x=23 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5950 N$11899 N$11900 "Straight Waveguide" sch_x=23 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5951 N$11901 N$11902 "Straight Waveguide" sch_x=23 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5952 N$11903 N$11904 "Straight Waveguide" sch_x=23 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5953 N$11905 N$11906 "Straight Waveguide" sch_x=23 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5954 N$11907 N$11908 "Straight Waveguide" sch_x=23 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5955 N$11909 N$11910 "Straight Waveguide" sch_x=23 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5956 N$11911 N$11912 "Straight Waveguide" sch_x=23 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5957 N$11913 N$11914 "Straight Waveguide" sch_x=21 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5958 N$11915 N$11916 "Straight Waveguide" sch_x=21 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5959 N$11917 N$11918 "Straight Waveguide" sch_x=21 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5960 N$11919 N$11920 "Straight Waveguide" sch_x=21 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5961 N$11921 N$11922 "Straight Waveguide" sch_x=21 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5962 N$11923 N$11924 "Straight Waveguide" sch_x=21 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5963 N$11925 N$11926 "Straight Waveguide" sch_x=19 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5964 N$11927 N$11928 "Straight Waveguide" sch_x=19 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5965 N$11929 N$11930 "Straight Waveguide" sch_x=19 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5966 N$11931 N$11932 "Straight Waveguide" sch_x=19 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5967 N$11933 N$11934 "Straight Waveguide" sch_x=17 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5968 N$11935 N$11936 "Straight Waveguide" sch_x=17 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5969 N$11938 N$11937 "Straight Waveguide" sch_x=21 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5970 N$11940 N$11939 "Straight Waveguide" sch_x=20 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5971 N$11942 N$11941 "Straight Waveguide" sch_x=19 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5972 N$11944 N$11943 "Straight Waveguide" sch_x=18 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5973 N$11946 N$11945 "Straight Waveguide" sch_x=17 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5974 N$11948 N$11947 "Straight Waveguide" sch_x=16 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5975 N$11950 N$11949 "Straight Waveguide" sch_x=15 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5976 N$11952 N$11951 "Straight Waveguide" sch_x=15 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5977 N$11954 N$11953 "Straight Waveguide" sch_x=16 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5978 N$11956 N$11955 "Straight Waveguide" sch_x=17 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5979 N$11958 N$11957 "Straight Waveguide" sch_x=18 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5980 N$11960 N$11959 "Straight Waveguide" sch_x=19 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5981 N$11962 N$11961 "Straight Waveguide" sch_x=20 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5982 N$11964 N$11963 "Straight Waveguide" sch_x=21 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5983 N$11966 N$11965 "Straight Waveguide" sch_x=22 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5984 N$11968 N$11967 "Straight Waveguide" sch_x=22 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5985 N$11969 N$11970 "Straight Waveguide" sch_x=-4 sch_y=-48.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5986 N$11971 N$11972 "Straight Waveguide" sch_x=-5 sch_y=-49.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5987 N$11973 N$11974 "Straight Waveguide" sch_x=-5 sch_y=-50.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5988 N$11975 N$11976 "Straight Waveguide" sch_x=-3 sch_y=-49.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5989 N$11977 N$11978 "Straight Waveguide" sch_x=-3 sch_y=-50.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5990 N$11979 N$11980 "Straight Waveguide" sch_x=-4 sch_y=-51.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5991 N$11981 N$11982 "Straight Waveguide" sch_x=0 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5992 N$11983 N$11984 "Straight Waveguide" sch_x=-1 sch_y=-48.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5993 N$11985 N$11986 "Straight Waveguide" sch_x=-1 sch_y=-49.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5994 N$11987 N$11988 "Straight Waveguide" sch_x=1 sch_y=-49.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5995 N$11989 N$11990 "Straight Waveguide" sch_x=1 sch_y=-48.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5996 N$11991 N$11992 "Straight Waveguide" sch_x=0 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5997 N$11993 N$11994 "Straight Waveguide" sch_x=0 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5998 N$11995 N$11996 "Straight Waveguide" sch_x=-1 sch_y=-50.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5999 N$11997 N$11998 "Straight Waveguide" sch_x=-1 sch_y=-51.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6000 N$11999 N$12000 "Straight Waveguide" sch_x=1 sch_y=-51.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6001 N$12001 N$12002 "Straight Waveguide" sch_x=1 sch_y=-50.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6002 N$12003 N$12004 "Straight Waveguide" sch_x=0 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6003 N$12005 N$12006 "Straight Waveguide" sch_x=4 sch_y=-48.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6004 N$12007 N$12008 "Straight Waveguide" sch_x=3 sch_y=-49.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6005 N$12009 N$12010 "Straight Waveguide" sch_x=3 sch_y=-50.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6006 N$12011 N$12012 "Straight Waveguide" sch_x=5 sch_y=-50.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6007 N$12013 N$12014 "Straight Waveguide" sch_x=5 sch_y=-49.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6008 N$12015 N$12016 "Straight Waveguide" sch_x=4 sch_y=-51.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6009 N$12017 N$12018 "Straight Waveguide" sch_x=-4 sch_y=-52.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6010 N$12019 N$12020 "Straight Waveguide" sch_x=-5 sch_y=-53.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6011 N$12021 N$12022 "Straight Waveguide" sch_x=-5 sch_y=-54.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6012 N$12023 N$12024 "Straight Waveguide" sch_x=-3 sch_y=-53.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6013 N$12025 N$12026 "Straight Waveguide" sch_x=-3 sch_y=-54.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6014 N$12027 N$12028 "Straight Waveguide" sch_x=-4 sch_y=-55.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6015 N$12029 N$12030 "Straight Waveguide" sch_x=0 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6016 N$12031 N$12032 "Straight Waveguide" sch_x=-1 sch_y=-52.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6017 N$12033 N$12034 "Straight Waveguide" sch_x=-1 sch_y=-53.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6018 N$12035 N$12036 "Straight Waveguide" sch_x=1 sch_y=-53.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6019 N$12037 N$12038 "Straight Waveguide" sch_x=1 sch_y=-52.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6020 N$12039 N$12040 "Straight Waveguide" sch_x=0 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6021 N$12041 N$12042 "Straight Waveguide" sch_x=0 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6022 N$12043 N$12044 "Straight Waveguide" sch_x=-1 sch_y=-54.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6023 N$12045 N$12046 "Straight Waveguide" sch_x=-1 sch_y=-55.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6024 N$12047 N$12048 "Straight Waveguide" sch_x=1 sch_y=-55.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6025 N$12049 N$12050 "Straight Waveguide" sch_x=1 sch_y=-54.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6026 N$12051 N$12052 "Straight Waveguide" sch_x=0 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6027 N$12053 N$12054 "Straight Waveguide" sch_x=4 sch_y=-52.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6028 N$12055 N$12056 "Straight Waveguide" sch_x=3 sch_y=-53.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6029 N$12057 N$12058 "Straight Waveguide" sch_x=3 sch_y=-54.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6030 N$12059 N$12060 "Straight Waveguide" sch_x=5 sch_y=-54.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6031 N$12061 N$12062 "Straight Waveguide" sch_x=5 sch_y=-53.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6032 N$12063 N$12064 "Straight Waveguide" sch_x=4 sch_y=-55.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6033 N$12066 N$12065 "Straight Waveguide" sch_x=-13 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6034 N$12068 N$12067 "Straight Waveguide" sch_x=-13 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6035 N$12070 N$12069 "Straight Waveguide" sch_x=-13 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6036 N$12072 N$12071 "Straight Waveguide" sch_x=-13 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6037 N$12074 N$12073 "Straight Waveguide" sch_x=-13 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6038 N$12076 N$12075 "Straight Waveguide" sch_x=-13 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6039 N$12078 N$12077 "Straight Waveguide" sch_x=-11 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6040 N$12080 N$12079 "Straight Waveguide" sch_x=-11 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6041 N$12082 N$12081 "Straight Waveguide" sch_x=-11 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6042 N$12084 N$12083 "Straight Waveguide" sch_x=-11 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6043 N$12086 N$12085 "Straight Waveguide" sch_x=-9 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6044 N$12088 N$12087 "Straight Waveguide" sch_x=-9 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6045 N$12089 N$12090 "Straight Waveguide" sch_x=-9 sch_y=-49.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6046 N$12091 N$12092 "Straight Waveguide" sch_x=-8 sch_y=-50.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6047 N$12093 N$12094 "Straight Waveguide" sch_x=-7 sch_y=-51.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6048 N$12095 N$12096 "Straight Waveguide" sch_x=-7 sch_y=-52.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6049 N$12097 N$12098 "Straight Waveguide" sch_x=-8 sch_y=-53.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6050 N$12099 N$12100 "Straight Waveguide" sch_x=-9 sch_y=-54.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6051 N$12101 N$12102 "Straight Waveguide" sch_x=-10 sch_y=-49.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6052 N$12103 N$12104 "Straight Waveguide" sch_x=-10 sch_y=-54.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6053 N$12105 N$12106 "Straight Waveguide" sch_x=13 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6054 N$12107 N$12108 "Straight Waveguide" sch_x=13 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6055 N$12109 N$12110 "Straight Waveguide" sch_x=13 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6056 N$12111 N$12112 "Straight Waveguide" sch_x=13 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6057 N$12113 N$12114 "Straight Waveguide" sch_x=13 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6058 N$12115 N$12116 "Straight Waveguide" sch_x=13 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6059 N$12117 N$12118 "Straight Waveguide" sch_x=11 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6060 N$12119 N$12120 "Straight Waveguide" sch_x=11 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6061 N$12121 N$12122 "Straight Waveguide" sch_x=11 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6062 N$12123 N$12124 "Straight Waveguide" sch_x=11 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6063 N$12125 N$12126 "Straight Waveguide" sch_x=9 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6064 N$12127 N$12128 "Straight Waveguide" sch_x=9 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6065 N$12130 N$12129 "Straight Waveguide" sch_x=9 sch_y=-49.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6066 N$12132 N$12131 "Straight Waveguide" sch_x=8 sch_y=-50.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6067 N$12134 N$12133 "Straight Waveguide" sch_x=7 sch_y=-51.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6068 N$12136 N$12135 "Straight Waveguide" sch_x=7 sch_y=-52.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6069 N$12138 N$12137 "Straight Waveguide" sch_x=8 sch_y=-53.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6070 N$12140 N$12139 "Straight Waveguide" sch_x=9 sch_y=-54.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6071 N$12142 N$12141 "Straight Waveguide" sch_x=10 sch_y=-49.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6072 N$12144 N$12143 "Straight Waveguide" sch_x=10 sch_y=-54.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6073 N$12145 N$12146 "Straight Waveguide" sch_x=-4 sch_y=-56.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6074 N$12147 N$12148 "Straight Waveguide" sch_x=-5 sch_y=-57.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6075 N$12149 N$12150 "Straight Waveguide" sch_x=-5 sch_y=-58.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6076 N$12151 N$12152 "Straight Waveguide" sch_x=-3 sch_y=-57.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6077 N$12153 N$12154 "Straight Waveguide" sch_x=-3 sch_y=-58.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6078 N$12155 N$12156 "Straight Waveguide" sch_x=-4 sch_y=-59.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6079 N$12157 N$12158 "Straight Waveguide" sch_x=0 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6080 N$12159 N$12160 "Straight Waveguide" sch_x=-1 sch_y=-56.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6081 N$12161 N$12162 "Straight Waveguide" sch_x=-1 sch_y=-57.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6082 N$12163 N$12164 "Straight Waveguide" sch_x=1 sch_y=-57.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6083 N$12165 N$12166 "Straight Waveguide" sch_x=1 sch_y=-56.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6084 N$12167 N$12168 "Straight Waveguide" sch_x=0 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6085 N$12169 N$12170 "Straight Waveguide" sch_x=0 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6086 N$12171 N$12172 "Straight Waveguide" sch_x=-1 sch_y=-58.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6087 N$12173 N$12174 "Straight Waveguide" sch_x=-1 sch_y=-59.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6088 N$12175 N$12176 "Straight Waveguide" sch_x=1 sch_y=-59.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6089 N$12177 N$12178 "Straight Waveguide" sch_x=1 sch_y=-58.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6090 N$12179 N$12180 "Straight Waveguide" sch_x=0 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6091 N$12181 N$12182 "Straight Waveguide" sch_x=4 sch_y=-56.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6092 N$12183 N$12184 "Straight Waveguide" sch_x=3 sch_y=-57.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6093 N$12185 N$12186 "Straight Waveguide" sch_x=3 sch_y=-58.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6094 N$12187 N$12188 "Straight Waveguide" sch_x=5 sch_y=-58.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6095 N$12189 N$12190 "Straight Waveguide" sch_x=5 sch_y=-57.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6096 N$12191 N$12192 "Straight Waveguide" sch_x=4 sch_y=-59.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6097 N$12193 N$12194 "Straight Waveguide" sch_x=-4 sch_y=-60.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6098 N$12195 N$12196 "Straight Waveguide" sch_x=-5 sch_y=-61.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6099 N$12197 N$12198 "Straight Waveguide" sch_x=-5 sch_y=-62.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6100 N$12199 N$12200 "Straight Waveguide" sch_x=-3 sch_y=-61.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6101 N$12201 N$12202 "Straight Waveguide" sch_x=-3 sch_y=-62.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6102 N$12203 N$12204 "Straight Waveguide" sch_x=-4 sch_y=-63.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6103 N$12205 N$12206 "Straight Waveguide" sch_x=0 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6104 N$12207 N$12208 "Straight Waveguide" sch_x=-1 sch_y=-60.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6105 N$12209 N$12210 "Straight Waveguide" sch_x=-1 sch_y=-61.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6106 N$12211 N$12212 "Straight Waveguide" sch_x=1 sch_y=-61.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6107 N$12213 N$12214 "Straight Waveguide" sch_x=1 sch_y=-60.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6108 N$12215 N$12216 "Straight Waveguide" sch_x=0 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6109 N$12217 N$12218 "Straight Waveguide" sch_x=0 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6110 N$12219 N$12220 "Straight Waveguide" sch_x=-1 sch_y=-62.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6111 N$12221 N$12222 "Straight Waveguide" sch_x=-1 sch_y=-63.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6112 N$12223 N$12224 "Straight Waveguide" sch_x=1 sch_y=-63.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6113 N$12225 N$12226 "Straight Waveguide" sch_x=1 sch_y=-62.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6114 N$12227 N$12228 "Straight Waveguide" sch_x=0 sch_y=-63.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6115 N$12229 N$12230 "Straight Waveguide" sch_x=4 sch_y=-60.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6116 N$12231 N$12232 "Straight Waveguide" sch_x=3 sch_y=-61.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6117 N$12233 N$12234 "Straight Waveguide" sch_x=3 sch_y=-62.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6118 N$12235 N$12236 "Straight Waveguide" sch_x=5 sch_y=-62.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6119 N$12237 N$12238 "Straight Waveguide" sch_x=5 sch_y=-61.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6120 N$12239 N$12240 "Straight Waveguide" sch_x=4 sch_y=-63.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6121 N$12242 N$12241 "Straight Waveguide" sch_x=-13 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6122 N$12244 N$12243 "Straight Waveguide" sch_x=-13 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6123 N$12246 N$12245 "Straight Waveguide" sch_x=-13 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6124 N$12248 N$12247 "Straight Waveguide" sch_x=-13 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6125 N$12250 N$12249 "Straight Waveguide" sch_x=-13 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6126 N$12252 N$12251 "Straight Waveguide" sch_x=-13 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6127 N$12254 N$12253 "Straight Waveguide" sch_x=-11 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6128 N$12256 N$12255 "Straight Waveguide" sch_x=-11 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6129 N$12258 N$12257 "Straight Waveguide" sch_x=-11 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6130 N$12260 N$12259 "Straight Waveguide" sch_x=-11 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6131 N$12262 N$12261 "Straight Waveguide" sch_x=-9 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6132 N$12264 N$12263 "Straight Waveguide" sch_x=-9 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6133 N$12265 N$12266 "Straight Waveguide" sch_x=-9 sch_y=-57.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6134 N$12267 N$12268 "Straight Waveguide" sch_x=-8 sch_y=-58.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6135 N$12269 N$12270 "Straight Waveguide" sch_x=-7 sch_y=-59.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6136 N$12271 N$12272 "Straight Waveguide" sch_x=-7 sch_y=-60.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6137 N$12273 N$12274 "Straight Waveguide" sch_x=-8 sch_y=-61.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6138 N$12275 N$12276 "Straight Waveguide" sch_x=-9 sch_y=-62.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6139 N$12277 N$12278 "Straight Waveguide" sch_x=-10 sch_y=-57.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6140 N$12279 N$12280 "Straight Waveguide" sch_x=-10 sch_y=-62.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6141 N$12281 N$12282 "Straight Waveguide" sch_x=13 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6142 N$12283 N$12284 "Straight Waveguide" sch_x=13 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6143 N$12285 N$12286 "Straight Waveguide" sch_x=13 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6144 N$12287 N$12288 "Straight Waveguide" sch_x=13 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6145 N$12289 N$12290 "Straight Waveguide" sch_x=13 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6146 N$12291 N$12292 "Straight Waveguide" sch_x=13 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6147 N$12293 N$12294 "Straight Waveguide" sch_x=11 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6148 N$12295 N$12296 "Straight Waveguide" sch_x=11 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6149 N$12297 N$12298 "Straight Waveguide" sch_x=11 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6150 N$12299 N$12300 "Straight Waveguide" sch_x=11 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6151 N$12301 N$12302 "Straight Waveguide" sch_x=9 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6152 N$12303 N$12304 "Straight Waveguide" sch_x=9 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6153 N$12306 N$12305 "Straight Waveguide" sch_x=9 sch_y=-57.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6154 N$12308 N$12307 "Straight Waveguide" sch_x=8 sch_y=-58.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6155 N$12310 N$12309 "Straight Waveguide" sch_x=7 sch_y=-59.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6156 N$12312 N$12311 "Straight Waveguide" sch_x=7 sch_y=-60.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6157 N$12314 N$12313 "Straight Waveguide" sch_x=8 sch_y=-61.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6158 N$12316 N$12315 "Straight Waveguide" sch_x=9 sch_y=-62.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6159 N$12318 N$12317 "Straight Waveguide" sch_x=10 sch_y=-57.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6160 N$12320 N$12319 "Straight Waveguide" sch_x=10 sch_y=-62.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6161 N$12322 N$12321 "Straight Waveguide" sch_x=-29 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6162 N$12324 N$12323 "Straight Waveguide" sch_x=-29 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6163 N$12326 N$12325 "Straight Waveguide" sch_x=-29 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6164 N$12328 N$12327 "Straight Waveguide" sch_x=-29 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6165 N$12330 N$12329 "Straight Waveguide" sch_x=-29 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6166 N$12332 N$12331 "Straight Waveguide" sch_x=-29 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6167 N$12334 N$12333 "Straight Waveguide" sch_x=-29 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6168 N$12336 N$12335 "Straight Waveguide" sch_x=-29 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6169 N$12338 N$12337 "Straight Waveguide" sch_x=-29 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6170 N$12340 N$12339 "Straight Waveguide" sch_x=-29 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6171 N$12342 N$12341 "Straight Waveguide" sch_x=-29 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6172 N$12344 N$12343 "Straight Waveguide" sch_x=-29 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6173 N$12346 N$12345 "Straight Waveguide" sch_x=-29 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6174 N$12348 N$12347 "Straight Waveguide" sch_x=-29 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6175 N$12350 N$12349 "Straight Waveguide" sch_x=-27 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6176 N$12352 N$12351 "Straight Waveguide" sch_x=-27 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6177 N$12354 N$12353 "Straight Waveguide" sch_x=-27 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6178 N$12356 N$12355 "Straight Waveguide" sch_x=-27 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6179 N$12358 N$12357 "Straight Waveguide" sch_x=-27 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6180 N$12360 N$12359 "Straight Waveguide" sch_x=-27 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6181 N$12362 N$12361 "Straight Waveguide" sch_x=-27 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6182 N$12364 N$12363 "Straight Waveguide" sch_x=-27 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6183 N$12366 N$12365 "Straight Waveguide" sch_x=-27 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6184 N$12368 N$12367 "Straight Waveguide" sch_x=-27 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6185 N$12370 N$12369 "Straight Waveguide" sch_x=-27 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6186 N$12372 N$12371 "Straight Waveguide" sch_x=-27 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6187 N$12374 N$12373 "Straight Waveguide" sch_x=-25 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6188 N$12376 N$12375 "Straight Waveguide" sch_x=-25 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6189 N$12378 N$12377 "Straight Waveguide" sch_x=-25 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6190 N$12380 N$12379 "Straight Waveguide" sch_x=-25 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6191 N$12382 N$12381 "Straight Waveguide" sch_x=-25 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6192 N$12384 N$12383 "Straight Waveguide" sch_x=-25 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6193 N$12386 N$12385 "Straight Waveguide" sch_x=-25 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6194 N$12388 N$12387 "Straight Waveguide" sch_x=-25 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6195 N$12390 N$12389 "Straight Waveguide" sch_x=-25 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6196 N$12392 N$12391 "Straight Waveguide" sch_x=-25 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6197 N$12394 N$12393 "Straight Waveguide" sch_x=-23 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6198 N$12396 N$12395 "Straight Waveguide" sch_x=-23 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6199 N$12398 N$12397 "Straight Waveguide" sch_x=-23 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6200 N$12400 N$12399 "Straight Waveguide" sch_x=-23 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6201 N$12402 N$12401 "Straight Waveguide" sch_x=-23 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6202 N$12404 N$12403 "Straight Waveguide" sch_x=-23 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6203 N$12406 N$12405 "Straight Waveguide" sch_x=-23 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6204 N$12408 N$12407 "Straight Waveguide" sch_x=-23 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6205 N$12410 N$12409 "Straight Waveguide" sch_x=-21 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6206 N$12412 N$12411 "Straight Waveguide" sch_x=-21 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6207 N$12414 N$12413 "Straight Waveguide" sch_x=-21 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6208 N$12416 N$12415 "Straight Waveguide" sch_x=-21 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6209 N$12418 N$12417 "Straight Waveguide" sch_x=-21 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6210 N$12420 N$12419 "Straight Waveguide" sch_x=-21 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6211 N$12422 N$12421 "Straight Waveguide" sch_x=-19 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6212 N$12424 N$12423 "Straight Waveguide" sch_x=-19 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6213 N$12426 N$12425 "Straight Waveguide" sch_x=-19 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6214 N$12428 N$12427 "Straight Waveguide" sch_x=-19 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6215 N$12430 N$12429 "Straight Waveguide" sch_x=-17 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6216 N$12432 N$12431 "Straight Waveguide" sch_x=-17 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6217 N$12433 N$12434 "Straight Waveguide" sch_x=-21 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6218 N$12435 N$12436 "Straight Waveguide" sch_x=-20 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6219 N$12437 N$12438 "Straight Waveguide" sch_x=-19 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6220 N$12439 N$12440 "Straight Waveguide" sch_x=-18 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6221 N$12441 N$12442 "Straight Waveguide" sch_x=-17 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6222 N$12443 N$12444 "Straight Waveguide" sch_x=-16 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6223 N$12445 N$12446 "Straight Waveguide" sch_x=-15 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6224 N$12447 N$12448 "Straight Waveguide" sch_x=-15 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6225 N$12449 N$12450 "Straight Waveguide" sch_x=-16 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6226 N$12451 N$12452 "Straight Waveguide" sch_x=-17 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6227 N$12453 N$12454 "Straight Waveguide" sch_x=-18 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6228 N$12455 N$12456 "Straight Waveguide" sch_x=-19 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6229 N$12457 N$12458 "Straight Waveguide" sch_x=-20 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6230 N$12459 N$12460 "Straight Waveguide" sch_x=-21 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6231 N$12461 N$12462 "Straight Waveguide" sch_x=-22 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6232 N$12463 N$12464 "Straight Waveguide" sch_x=-22 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6233 N$12465 N$12466 "Straight Waveguide" sch_x=29 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6234 N$12467 N$12468 "Straight Waveguide" sch_x=29 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6235 N$12469 N$12470 "Straight Waveguide" sch_x=29 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6236 N$12471 N$12472 "Straight Waveguide" sch_x=29 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6237 N$12473 N$12474 "Straight Waveguide" sch_x=29 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6238 N$12475 N$12476 "Straight Waveguide" sch_x=29 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6239 N$12477 N$12478 "Straight Waveguide" sch_x=29 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6240 N$12479 N$12480 "Straight Waveguide" sch_x=29 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6241 N$12481 N$12482 "Straight Waveguide" sch_x=29 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6242 N$12483 N$12484 "Straight Waveguide" sch_x=29 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6243 N$12485 N$12486 "Straight Waveguide" sch_x=29 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6244 N$12487 N$12488 "Straight Waveguide" sch_x=29 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6245 N$12489 N$12490 "Straight Waveguide" sch_x=29 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6246 N$12491 N$12492 "Straight Waveguide" sch_x=29 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6247 N$12493 N$12494 "Straight Waveguide" sch_x=27 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6248 N$12495 N$12496 "Straight Waveguide" sch_x=27 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6249 N$12497 N$12498 "Straight Waveguide" sch_x=27 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6250 N$12499 N$12500 "Straight Waveguide" sch_x=27 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6251 N$12501 N$12502 "Straight Waveguide" sch_x=27 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6252 N$12503 N$12504 "Straight Waveguide" sch_x=27 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6253 N$12505 N$12506 "Straight Waveguide" sch_x=27 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6254 N$12507 N$12508 "Straight Waveguide" sch_x=27 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6255 N$12509 N$12510 "Straight Waveguide" sch_x=27 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6256 N$12511 N$12512 "Straight Waveguide" sch_x=27 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6257 N$12513 N$12514 "Straight Waveguide" sch_x=27 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6258 N$12515 N$12516 "Straight Waveguide" sch_x=27 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6259 N$12517 N$12518 "Straight Waveguide" sch_x=25 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6260 N$12519 N$12520 "Straight Waveguide" sch_x=25 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6261 N$12521 N$12522 "Straight Waveguide" sch_x=25 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6262 N$12523 N$12524 "Straight Waveguide" sch_x=25 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6263 N$12525 N$12526 "Straight Waveguide" sch_x=25 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6264 N$12527 N$12528 "Straight Waveguide" sch_x=25 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6265 N$12529 N$12530 "Straight Waveguide" sch_x=25 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6266 N$12531 N$12532 "Straight Waveguide" sch_x=25 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6267 N$12533 N$12534 "Straight Waveguide" sch_x=25 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6268 N$12535 N$12536 "Straight Waveguide" sch_x=25 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6269 N$12537 N$12538 "Straight Waveguide" sch_x=23 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6270 N$12539 N$12540 "Straight Waveguide" sch_x=23 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6271 N$12541 N$12542 "Straight Waveguide" sch_x=23 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6272 N$12543 N$12544 "Straight Waveguide" sch_x=23 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6273 N$12545 N$12546 "Straight Waveguide" sch_x=23 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6274 N$12547 N$12548 "Straight Waveguide" sch_x=23 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6275 N$12549 N$12550 "Straight Waveguide" sch_x=23 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6276 N$12551 N$12552 "Straight Waveguide" sch_x=23 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6277 N$12553 N$12554 "Straight Waveguide" sch_x=21 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6278 N$12555 N$12556 "Straight Waveguide" sch_x=21 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6279 N$12557 N$12558 "Straight Waveguide" sch_x=21 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6280 N$12559 N$12560 "Straight Waveguide" sch_x=21 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6281 N$12561 N$12562 "Straight Waveguide" sch_x=21 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6282 N$12563 N$12564 "Straight Waveguide" sch_x=21 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6283 N$12565 N$12566 "Straight Waveguide" sch_x=19 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6284 N$12567 N$12568 "Straight Waveguide" sch_x=19 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6285 N$12569 N$12570 "Straight Waveguide" sch_x=19 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6286 N$12571 N$12572 "Straight Waveguide" sch_x=19 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6287 N$12573 N$12574 "Straight Waveguide" sch_x=17 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6288 N$12575 N$12576 "Straight Waveguide" sch_x=17 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6289 N$12578 N$12577 "Straight Waveguide" sch_x=21 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6290 N$12580 N$12579 "Straight Waveguide" sch_x=20 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6291 N$12582 N$12581 "Straight Waveguide" sch_x=19 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6292 N$12584 N$12583 "Straight Waveguide" sch_x=18 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6293 N$12586 N$12585 "Straight Waveguide" sch_x=17 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6294 N$12588 N$12587 "Straight Waveguide" sch_x=16 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6295 N$12590 N$12589 "Straight Waveguide" sch_x=15 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6296 N$12592 N$12591 "Straight Waveguide" sch_x=15 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6297 N$12594 N$12593 "Straight Waveguide" sch_x=16 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6298 N$12596 N$12595 "Straight Waveguide" sch_x=17 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6299 N$12598 N$12597 "Straight Waveguide" sch_x=18 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6300 N$12600 N$12599 "Straight Waveguide" sch_x=19 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6301 N$12602 N$12601 "Straight Waveguide" sch_x=20 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6302 N$12604 N$12603 "Straight Waveguide" sch_x=21 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6303 N$12606 N$12605 "Straight Waveguide" sch_x=22 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6304 N$12608 N$12607 "Straight Waveguide" sch_x=22 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6305 N$12610 N$12609 "Straight Waveguide" sch_x=-61 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6306 N$12612 N$12611 "Straight Waveguide" sch_x=-61 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6307 N$12614 N$12613 "Straight Waveguide" sch_x=-61 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6308 N$12616 N$12615 "Straight Waveguide" sch_x=-61 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6309 N$12618 N$12617 "Straight Waveguide" sch_x=-61 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6310 N$12620 N$12619 "Straight Waveguide" sch_x=-61 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6311 N$12622 N$12621 "Straight Waveguide" sch_x=-61 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6312 N$12624 N$12623 "Straight Waveguide" sch_x=-61 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6313 N$12626 N$12625 "Straight Waveguide" sch_x=-61 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6314 N$12628 N$12627 "Straight Waveguide" sch_x=-61 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6315 N$12630 N$12629 "Straight Waveguide" sch_x=-61 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6316 N$12632 N$12631 "Straight Waveguide" sch_x=-61 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6317 N$12634 N$12633 "Straight Waveguide" sch_x=-61 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6318 N$12636 N$12635 "Straight Waveguide" sch_x=-61 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6319 N$12638 N$12637 "Straight Waveguide" sch_x=-61 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6320 N$12640 N$12639 "Straight Waveguide" sch_x=-61 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6321 N$12642 N$12641 "Straight Waveguide" sch_x=-61 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6322 N$12644 N$12643 "Straight Waveguide" sch_x=-61 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6323 N$12646 N$12645 "Straight Waveguide" sch_x=-61 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6324 N$12648 N$12647 "Straight Waveguide" sch_x=-61 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6325 N$12650 N$12649 "Straight Waveguide" sch_x=-61 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6326 N$12652 N$12651 "Straight Waveguide" sch_x=-61 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6327 N$12654 N$12653 "Straight Waveguide" sch_x=-61 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6328 N$12656 N$12655 "Straight Waveguide" sch_x=-61 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6329 N$12658 N$12657 "Straight Waveguide" sch_x=-61 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6330 N$12660 N$12659 "Straight Waveguide" sch_x=-61 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6331 N$12662 N$12661 "Straight Waveguide" sch_x=-61 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6332 N$12664 N$12663 "Straight Waveguide" sch_x=-61 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6333 N$12666 N$12665 "Straight Waveguide" sch_x=-61 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6334 N$12668 N$12667 "Straight Waveguide" sch_x=-61 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6335 N$12670 N$12669 "Straight Waveguide" sch_x=-59 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6336 N$12672 N$12671 "Straight Waveguide" sch_x=-59 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6337 N$12674 N$12673 "Straight Waveguide" sch_x=-59 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6338 N$12676 N$12675 "Straight Waveguide" sch_x=-59 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6339 N$12678 N$12677 "Straight Waveguide" sch_x=-59 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6340 N$12680 N$12679 "Straight Waveguide" sch_x=-59 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6341 N$12682 N$12681 "Straight Waveguide" sch_x=-59 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6342 N$12684 N$12683 "Straight Waveguide" sch_x=-59 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6343 N$12686 N$12685 "Straight Waveguide" sch_x=-59 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6344 N$12688 N$12687 "Straight Waveguide" sch_x=-59 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6345 N$12690 N$12689 "Straight Waveguide" sch_x=-59 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6346 N$12692 N$12691 "Straight Waveguide" sch_x=-59 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6347 N$12694 N$12693 "Straight Waveguide" sch_x=-59 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6348 N$12696 N$12695 "Straight Waveguide" sch_x=-59 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6349 N$12698 N$12697 "Straight Waveguide" sch_x=-59 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6350 N$12700 N$12699 "Straight Waveguide" sch_x=-59 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6351 N$12702 N$12701 "Straight Waveguide" sch_x=-59 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6352 N$12704 N$12703 "Straight Waveguide" sch_x=-59 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6353 N$12706 N$12705 "Straight Waveguide" sch_x=-59 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6354 N$12708 N$12707 "Straight Waveguide" sch_x=-59 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6355 N$12710 N$12709 "Straight Waveguide" sch_x=-59 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6356 N$12712 N$12711 "Straight Waveguide" sch_x=-59 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6357 N$12714 N$12713 "Straight Waveguide" sch_x=-59 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6358 N$12716 N$12715 "Straight Waveguide" sch_x=-59 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6359 N$12718 N$12717 "Straight Waveguide" sch_x=-59 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6360 N$12720 N$12719 "Straight Waveguide" sch_x=-59 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6361 N$12722 N$12721 "Straight Waveguide" sch_x=-59 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6362 N$12724 N$12723 "Straight Waveguide" sch_x=-59 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6363 N$12726 N$12725 "Straight Waveguide" sch_x=-57 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6364 N$12728 N$12727 "Straight Waveguide" sch_x=-57 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6365 N$12730 N$12729 "Straight Waveguide" sch_x=-57 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6366 N$12732 N$12731 "Straight Waveguide" sch_x=-57 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6367 N$12734 N$12733 "Straight Waveguide" sch_x=-57 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6368 N$12736 N$12735 "Straight Waveguide" sch_x=-57 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6369 N$12738 N$12737 "Straight Waveguide" sch_x=-57 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6370 N$12740 N$12739 "Straight Waveguide" sch_x=-57 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6371 N$12742 N$12741 "Straight Waveguide" sch_x=-57 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6372 N$12744 N$12743 "Straight Waveguide" sch_x=-57 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6373 N$12746 N$12745 "Straight Waveguide" sch_x=-57 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6374 N$12748 N$12747 "Straight Waveguide" sch_x=-57 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6375 N$12750 N$12749 "Straight Waveguide" sch_x=-57 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6376 N$12752 N$12751 "Straight Waveguide" sch_x=-57 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6377 N$12754 N$12753 "Straight Waveguide" sch_x=-57 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6378 N$12756 N$12755 "Straight Waveguide" sch_x=-57 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6379 N$12758 N$12757 "Straight Waveguide" sch_x=-57 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6380 N$12760 N$12759 "Straight Waveguide" sch_x=-57 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6381 N$12762 N$12761 "Straight Waveguide" sch_x=-57 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6382 N$12764 N$12763 "Straight Waveguide" sch_x=-57 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6383 N$12766 N$12765 "Straight Waveguide" sch_x=-57 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6384 N$12768 N$12767 "Straight Waveguide" sch_x=-57 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6385 N$12770 N$12769 "Straight Waveguide" sch_x=-57 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6386 N$12772 N$12771 "Straight Waveguide" sch_x=-57 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6387 N$12774 N$12773 "Straight Waveguide" sch_x=-57 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6388 N$12776 N$12775 "Straight Waveguide" sch_x=-57 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6389 N$12778 N$12777 "Straight Waveguide" sch_x=-55 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6390 N$12780 N$12779 "Straight Waveguide" sch_x=-55 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6391 N$12782 N$12781 "Straight Waveguide" sch_x=-55 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6392 N$12784 N$12783 "Straight Waveguide" sch_x=-55 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6393 N$12786 N$12785 "Straight Waveguide" sch_x=-55 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6394 N$12788 N$12787 "Straight Waveguide" sch_x=-55 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6395 N$12790 N$12789 "Straight Waveguide" sch_x=-55 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6396 N$12792 N$12791 "Straight Waveguide" sch_x=-55 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6397 N$12794 N$12793 "Straight Waveguide" sch_x=-55 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6398 N$12796 N$12795 "Straight Waveguide" sch_x=-55 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6399 N$12798 N$12797 "Straight Waveguide" sch_x=-55 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6400 N$12800 N$12799 "Straight Waveguide" sch_x=-55 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6401 N$12802 N$12801 "Straight Waveguide" sch_x=-55 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6402 N$12804 N$12803 "Straight Waveguide" sch_x=-55 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6403 N$12806 N$12805 "Straight Waveguide" sch_x=-55 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6404 N$12808 N$12807 "Straight Waveguide" sch_x=-55 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6405 N$12810 N$12809 "Straight Waveguide" sch_x=-55 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6406 N$12812 N$12811 "Straight Waveguide" sch_x=-55 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6407 N$12814 N$12813 "Straight Waveguide" sch_x=-55 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6408 N$12816 N$12815 "Straight Waveguide" sch_x=-55 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6409 N$12818 N$12817 "Straight Waveguide" sch_x=-55 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6410 N$12820 N$12819 "Straight Waveguide" sch_x=-55 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6411 N$12822 N$12821 "Straight Waveguide" sch_x=-55 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6412 N$12824 N$12823 "Straight Waveguide" sch_x=-55 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6413 N$12826 N$12825 "Straight Waveguide" sch_x=-53 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6414 N$12828 N$12827 "Straight Waveguide" sch_x=-53 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6415 N$12830 N$12829 "Straight Waveguide" sch_x=-53 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6416 N$12832 N$12831 "Straight Waveguide" sch_x=-53 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6417 N$12834 N$12833 "Straight Waveguide" sch_x=-53 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6418 N$12836 N$12835 "Straight Waveguide" sch_x=-53 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6419 N$12838 N$12837 "Straight Waveguide" sch_x=-53 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6420 N$12840 N$12839 "Straight Waveguide" sch_x=-53 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6421 N$12842 N$12841 "Straight Waveguide" sch_x=-53 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6422 N$12844 N$12843 "Straight Waveguide" sch_x=-53 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6423 N$12846 N$12845 "Straight Waveguide" sch_x=-53 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6424 N$12848 N$12847 "Straight Waveguide" sch_x=-53 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6425 N$12850 N$12849 "Straight Waveguide" sch_x=-53 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6426 N$12852 N$12851 "Straight Waveguide" sch_x=-53 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6427 N$12854 N$12853 "Straight Waveguide" sch_x=-53 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6428 N$12856 N$12855 "Straight Waveguide" sch_x=-53 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6429 N$12858 N$12857 "Straight Waveguide" sch_x=-53 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6430 N$12860 N$12859 "Straight Waveguide" sch_x=-53 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6431 N$12862 N$12861 "Straight Waveguide" sch_x=-53 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6432 N$12864 N$12863 "Straight Waveguide" sch_x=-53 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6433 N$12866 N$12865 "Straight Waveguide" sch_x=-53 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6434 N$12868 N$12867 "Straight Waveguide" sch_x=-53 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6435 N$12870 N$12869 "Straight Waveguide" sch_x=-51 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6436 N$12872 N$12871 "Straight Waveguide" sch_x=-51 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6437 N$12874 N$12873 "Straight Waveguide" sch_x=-51 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6438 N$12876 N$12875 "Straight Waveguide" sch_x=-51 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6439 N$12878 N$12877 "Straight Waveguide" sch_x=-51 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6440 N$12880 N$12879 "Straight Waveguide" sch_x=-51 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6441 N$12882 N$12881 "Straight Waveguide" sch_x=-51 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6442 N$12884 N$12883 "Straight Waveguide" sch_x=-51 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6443 N$12886 N$12885 "Straight Waveguide" sch_x=-51 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6444 N$12888 N$12887 "Straight Waveguide" sch_x=-51 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6445 N$12890 N$12889 "Straight Waveguide" sch_x=-51 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6446 N$12892 N$12891 "Straight Waveguide" sch_x=-51 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6447 N$12894 N$12893 "Straight Waveguide" sch_x=-51 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6448 N$12896 N$12895 "Straight Waveguide" sch_x=-51 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6449 N$12898 N$12897 "Straight Waveguide" sch_x=-51 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6450 N$12900 N$12899 "Straight Waveguide" sch_x=-51 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6451 N$12902 N$12901 "Straight Waveguide" sch_x=-51 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6452 N$12904 N$12903 "Straight Waveguide" sch_x=-51 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6453 N$12906 N$12905 "Straight Waveguide" sch_x=-51 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6454 N$12908 N$12907 "Straight Waveguide" sch_x=-51 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6455 N$12910 N$12909 "Straight Waveguide" sch_x=-49 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6456 N$12912 N$12911 "Straight Waveguide" sch_x=-49 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6457 N$12914 N$12913 "Straight Waveguide" sch_x=-49 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6458 N$12916 N$12915 "Straight Waveguide" sch_x=-49 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6459 N$12918 N$12917 "Straight Waveguide" sch_x=-49 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6460 N$12920 N$12919 "Straight Waveguide" sch_x=-49 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6461 N$12922 N$12921 "Straight Waveguide" sch_x=-49 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6462 N$12924 N$12923 "Straight Waveguide" sch_x=-49 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6463 N$12926 N$12925 "Straight Waveguide" sch_x=-49 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6464 N$12928 N$12927 "Straight Waveguide" sch_x=-49 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6465 N$12930 N$12929 "Straight Waveguide" sch_x=-49 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6466 N$12932 N$12931 "Straight Waveguide" sch_x=-49 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6467 N$12934 N$12933 "Straight Waveguide" sch_x=-49 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6468 N$12936 N$12935 "Straight Waveguide" sch_x=-49 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6469 N$12938 N$12937 "Straight Waveguide" sch_x=-49 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6470 N$12940 N$12939 "Straight Waveguide" sch_x=-49 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6471 N$12942 N$12941 "Straight Waveguide" sch_x=-49 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6472 N$12944 N$12943 "Straight Waveguide" sch_x=-49 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6473 N$12946 N$12945 "Straight Waveguide" sch_x=-47 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6474 N$12948 N$12947 "Straight Waveguide" sch_x=-47 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6475 N$12950 N$12949 "Straight Waveguide" sch_x=-47 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6476 N$12952 N$12951 "Straight Waveguide" sch_x=-47 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6477 N$12954 N$12953 "Straight Waveguide" sch_x=-47 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6478 N$12956 N$12955 "Straight Waveguide" sch_x=-47 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6479 N$12958 N$12957 "Straight Waveguide" sch_x=-47 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6480 N$12960 N$12959 "Straight Waveguide" sch_x=-47 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6481 N$12962 N$12961 "Straight Waveguide" sch_x=-47 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6482 N$12964 N$12963 "Straight Waveguide" sch_x=-47 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6483 N$12966 N$12965 "Straight Waveguide" sch_x=-47 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6484 N$12968 N$12967 "Straight Waveguide" sch_x=-47 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6485 N$12970 N$12969 "Straight Waveguide" sch_x=-47 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6486 N$12972 N$12971 "Straight Waveguide" sch_x=-47 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6487 N$12974 N$12973 "Straight Waveguide" sch_x=-47 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6488 N$12976 N$12975 "Straight Waveguide" sch_x=-47 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6489 N$12978 N$12977 "Straight Waveguide" sch_x=-45 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6490 N$12980 N$12979 "Straight Waveguide" sch_x=-45 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6491 N$12982 N$12981 "Straight Waveguide" sch_x=-45 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6492 N$12984 N$12983 "Straight Waveguide" sch_x=-45 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6493 N$12986 N$12985 "Straight Waveguide" sch_x=-45 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6494 N$12988 N$12987 "Straight Waveguide" sch_x=-45 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6495 N$12990 N$12989 "Straight Waveguide" sch_x=-45 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6496 N$12992 N$12991 "Straight Waveguide" sch_x=-45 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6497 N$12994 N$12993 "Straight Waveguide" sch_x=-45 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6498 N$12996 N$12995 "Straight Waveguide" sch_x=-45 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6499 N$12998 N$12997 "Straight Waveguide" sch_x=-45 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6500 N$13000 N$12999 "Straight Waveguide" sch_x=-45 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6501 N$13002 N$13001 "Straight Waveguide" sch_x=-45 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6502 N$13004 N$13003 "Straight Waveguide" sch_x=-45 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6503 N$13006 N$13005 "Straight Waveguide" sch_x=-43 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6504 N$13008 N$13007 "Straight Waveguide" sch_x=-43 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6505 N$13010 N$13009 "Straight Waveguide" sch_x=-43 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6506 N$13012 N$13011 "Straight Waveguide" sch_x=-43 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6507 N$13014 N$13013 "Straight Waveguide" sch_x=-43 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6508 N$13016 N$13015 "Straight Waveguide" sch_x=-43 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6509 N$13018 N$13017 "Straight Waveguide" sch_x=-43 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6510 N$13020 N$13019 "Straight Waveguide" sch_x=-43 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6511 N$13022 N$13021 "Straight Waveguide" sch_x=-43 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6512 N$13024 N$13023 "Straight Waveguide" sch_x=-43 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6513 N$13026 N$13025 "Straight Waveguide" sch_x=-43 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6514 N$13028 N$13027 "Straight Waveguide" sch_x=-43 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6515 N$13030 N$13029 "Straight Waveguide" sch_x=-41 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6516 N$13032 N$13031 "Straight Waveguide" sch_x=-41 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6517 N$13034 N$13033 "Straight Waveguide" sch_x=-41 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6518 N$13036 N$13035 "Straight Waveguide" sch_x=-41 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6519 N$13038 N$13037 "Straight Waveguide" sch_x=-41 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6520 N$13040 N$13039 "Straight Waveguide" sch_x=-41 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6521 N$13042 N$13041 "Straight Waveguide" sch_x=-41 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6522 N$13044 N$13043 "Straight Waveguide" sch_x=-41 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6523 N$13046 N$13045 "Straight Waveguide" sch_x=-41 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6524 N$13048 N$13047 "Straight Waveguide" sch_x=-41 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6525 N$13050 N$13049 "Straight Waveguide" sch_x=-39 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6526 N$13052 N$13051 "Straight Waveguide" sch_x=-39 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6527 N$13054 N$13053 "Straight Waveguide" sch_x=-39 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6528 N$13056 N$13055 "Straight Waveguide" sch_x=-39 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6529 N$13058 N$13057 "Straight Waveguide" sch_x=-39 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6530 N$13060 N$13059 "Straight Waveguide" sch_x=-39 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6531 N$13062 N$13061 "Straight Waveguide" sch_x=-39 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6532 N$13064 N$13063 "Straight Waveguide" sch_x=-39 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6533 N$13066 N$13065 "Straight Waveguide" sch_x=-37 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6534 N$13068 N$13067 "Straight Waveguide" sch_x=-37 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6535 N$13070 N$13069 "Straight Waveguide" sch_x=-37 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6536 N$13072 N$13071 "Straight Waveguide" sch_x=-37 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6537 N$13074 N$13073 "Straight Waveguide" sch_x=-37 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6538 N$13076 N$13075 "Straight Waveguide" sch_x=-37 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6539 N$13078 N$13077 "Straight Waveguide" sch_x=-35 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6540 N$13080 N$13079 "Straight Waveguide" sch_x=-35 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6541 N$13082 N$13081 "Straight Waveguide" sch_x=-35 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6542 N$13084 N$13083 "Straight Waveguide" sch_x=-35 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6543 N$13086 N$13085 "Straight Waveguide" sch_x=-33 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6544 N$13088 N$13087 "Straight Waveguide" sch_x=-33 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6545 N$13089 N$13090 "Straight Waveguide" sch_x=-45 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6546 N$13091 N$13092 "Straight Waveguide" sch_x=-44 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6547 N$13093 N$13094 "Straight Waveguide" sch_x=-43 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6548 N$13095 N$13096 "Straight Waveguide" sch_x=-42 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6549 N$13097 N$13098 "Straight Waveguide" sch_x=-41 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6550 N$13099 N$13100 "Straight Waveguide" sch_x=-40 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6551 N$13101 N$13102 "Straight Waveguide" sch_x=-39 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6552 N$13103 N$13104 "Straight Waveguide" sch_x=-38 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6553 N$13105 N$13106 "Straight Waveguide" sch_x=-37 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6554 N$13107 N$13108 "Straight Waveguide" sch_x=-36 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6555 N$13109 N$13110 "Straight Waveguide" sch_x=-35 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6556 N$13111 N$13112 "Straight Waveguide" sch_x=-34 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6557 N$13113 N$13114 "Straight Waveguide" sch_x=-33 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6558 N$13115 N$13116 "Straight Waveguide" sch_x=-32 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6559 N$13117 N$13118 "Straight Waveguide" sch_x=-31 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6560 N$13119 N$13120 "Straight Waveguide" sch_x=-31 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6561 N$13121 N$13122 "Straight Waveguide" sch_x=-32 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6562 N$13123 N$13124 "Straight Waveguide" sch_x=-33 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6563 N$13125 N$13126 "Straight Waveguide" sch_x=-34 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6564 N$13127 N$13128 "Straight Waveguide" sch_x=-35 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6565 N$13129 N$13130 "Straight Waveguide" sch_x=-36 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6566 N$13131 N$13132 "Straight Waveguide" sch_x=-37 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6567 N$13133 N$13134 "Straight Waveguide" sch_x=-38 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6568 N$13135 N$13136 "Straight Waveguide" sch_x=-39 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6569 N$13137 N$13138 "Straight Waveguide" sch_x=-40 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6570 N$13139 N$13140 "Straight Waveguide" sch_x=-41 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6571 N$13141 N$13142 "Straight Waveguide" sch_x=-42 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6572 N$13143 N$13144 "Straight Waveguide" sch_x=-43 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6573 N$13145 N$13146 "Straight Waveguide" sch_x=-44 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6574 N$13147 N$13148 "Straight Waveguide" sch_x=-45 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6575 N$13149 N$13150 "Straight Waveguide" sch_x=-46 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6576 N$13151 N$13152 "Straight Waveguide" sch_x=-46 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6577 N$13153 N$13154 "Straight Waveguide" sch_x=61 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6578 N$13155 N$13156 "Straight Waveguide" sch_x=61 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6579 N$13157 N$13158 "Straight Waveguide" sch_x=61 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6580 N$13159 N$13160 "Straight Waveguide" sch_x=61 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6581 N$13161 N$13162 "Straight Waveguide" sch_x=61 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6582 N$13163 N$13164 "Straight Waveguide" sch_x=61 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6583 N$13165 N$13166 "Straight Waveguide" sch_x=61 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6584 N$13167 N$13168 "Straight Waveguide" sch_x=61 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6585 N$13169 N$13170 "Straight Waveguide" sch_x=61 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6586 N$13171 N$13172 "Straight Waveguide" sch_x=61 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6587 N$13173 N$13174 "Straight Waveguide" sch_x=61 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6588 N$13175 N$13176 "Straight Waveguide" sch_x=61 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6589 N$13177 N$13178 "Straight Waveguide" sch_x=61 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6590 N$13179 N$13180 "Straight Waveguide" sch_x=61 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6591 N$13181 N$13182 "Straight Waveguide" sch_x=61 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6592 N$13183 N$13184 "Straight Waveguide" sch_x=61 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6593 N$13185 N$13186 "Straight Waveguide" sch_x=61 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6594 N$13187 N$13188 "Straight Waveguide" sch_x=61 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6595 N$13189 N$13190 "Straight Waveguide" sch_x=61 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6596 N$13191 N$13192 "Straight Waveguide" sch_x=61 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6597 N$13193 N$13194 "Straight Waveguide" sch_x=61 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6598 N$13195 N$13196 "Straight Waveguide" sch_x=61 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6599 N$13197 N$13198 "Straight Waveguide" sch_x=61 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6600 N$13199 N$13200 "Straight Waveguide" sch_x=61 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6601 N$13201 N$13202 "Straight Waveguide" sch_x=61 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6602 N$13203 N$13204 "Straight Waveguide" sch_x=61 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6603 N$13205 N$13206 "Straight Waveguide" sch_x=61 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6604 N$13207 N$13208 "Straight Waveguide" sch_x=61 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6605 N$13209 N$13210 "Straight Waveguide" sch_x=61 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6606 N$13211 N$13212 "Straight Waveguide" sch_x=61 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6607 N$13213 N$13214 "Straight Waveguide" sch_x=59 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6608 N$13215 N$13216 "Straight Waveguide" sch_x=59 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6609 N$13217 N$13218 "Straight Waveguide" sch_x=59 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6610 N$13219 N$13220 "Straight Waveguide" sch_x=59 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6611 N$13221 N$13222 "Straight Waveguide" sch_x=59 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6612 N$13223 N$13224 "Straight Waveguide" sch_x=59 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6613 N$13225 N$13226 "Straight Waveguide" sch_x=59 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6614 N$13227 N$13228 "Straight Waveguide" sch_x=59 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6615 N$13229 N$13230 "Straight Waveguide" sch_x=59 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6616 N$13231 N$13232 "Straight Waveguide" sch_x=59 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6617 N$13233 N$13234 "Straight Waveguide" sch_x=59 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6618 N$13235 N$13236 "Straight Waveguide" sch_x=59 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6619 N$13237 N$13238 "Straight Waveguide" sch_x=59 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6620 N$13239 N$13240 "Straight Waveguide" sch_x=59 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6621 N$13241 N$13242 "Straight Waveguide" sch_x=59 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6622 N$13243 N$13244 "Straight Waveguide" sch_x=59 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6623 N$13245 N$13246 "Straight Waveguide" sch_x=59 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6624 N$13247 N$13248 "Straight Waveguide" sch_x=59 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6625 N$13249 N$13250 "Straight Waveguide" sch_x=59 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6626 N$13251 N$13252 "Straight Waveguide" sch_x=59 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6627 N$13253 N$13254 "Straight Waveguide" sch_x=59 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6628 N$13255 N$13256 "Straight Waveguide" sch_x=59 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6629 N$13257 N$13258 "Straight Waveguide" sch_x=59 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6630 N$13259 N$13260 "Straight Waveguide" sch_x=59 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6631 N$13261 N$13262 "Straight Waveguide" sch_x=59 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6632 N$13263 N$13264 "Straight Waveguide" sch_x=59 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6633 N$13265 N$13266 "Straight Waveguide" sch_x=59 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6634 N$13267 N$13268 "Straight Waveguide" sch_x=59 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6635 N$13269 N$13270 "Straight Waveguide" sch_x=57 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6636 N$13271 N$13272 "Straight Waveguide" sch_x=57 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6637 N$13273 N$13274 "Straight Waveguide" sch_x=57 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6638 N$13275 N$13276 "Straight Waveguide" sch_x=57 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6639 N$13277 N$13278 "Straight Waveguide" sch_x=57 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6640 N$13279 N$13280 "Straight Waveguide" sch_x=57 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6641 N$13281 N$13282 "Straight Waveguide" sch_x=57 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6642 N$13283 N$13284 "Straight Waveguide" sch_x=57 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6643 N$13285 N$13286 "Straight Waveguide" sch_x=57 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6644 N$13287 N$13288 "Straight Waveguide" sch_x=57 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6645 N$13289 N$13290 "Straight Waveguide" sch_x=57 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6646 N$13291 N$13292 "Straight Waveguide" sch_x=57 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6647 N$13293 N$13294 "Straight Waveguide" sch_x=57 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6648 N$13295 N$13296 "Straight Waveguide" sch_x=57 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6649 N$13297 N$13298 "Straight Waveguide" sch_x=57 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6650 N$13299 N$13300 "Straight Waveguide" sch_x=57 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6651 N$13301 N$13302 "Straight Waveguide" sch_x=57 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6652 N$13303 N$13304 "Straight Waveguide" sch_x=57 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6653 N$13305 N$13306 "Straight Waveguide" sch_x=57 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6654 N$13307 N$13308 "Straight Waveguide" sch_x=57 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6655 N$13309 N$13310 "Straight Waveguide" sch_x=57 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6656 N$13311 N$13312 "Straight Waveguide" sch_x=57 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6657 N$13313 N$13314 "Straight Waveguide" sch_x=57 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6658 N$13315 N$13316 "Straight Waveguide" sch_x=57 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6659 N$13317 N$13318 "Straight Waveguide" sch_x=57 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6660 N$13319 N$13320 "Straight Waveguide" sch_x=57 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6661 N$13321 N$13322 "Straight Waveguide" sch_x=55 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6662 N$13323 N$13324 "Straight Waveguide" sch_x=55 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6663 N$13325 N$13326 "Straight Waveguide" sch_x=55 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6664 N$13327 N$13328 "Straight Waveguide" sch_x=55 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6665 N$13329 N$13330 "Straight Waveguide" sch_x=55 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6666 N$13331 N$13332 "Straight Waveguide" sch_x=55 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6667 N$13333 N$13334 "Straight Waveguide" sch_x=55 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6668 N$13335 N$13336 "Straight Waveguide" sch_x=55 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6669 N$13337 N$13338 "Straight Waveguide" sch_x=55 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6670 N$13339 N$13340 "Straight Waveguide" sch_x=55 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6671 N$13341 N$13342 "Straight Waveguide" sch_x=55 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6672 N$13343 N$13344 "Straight Waveguide" sch_x=55 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6673 N$13345 N$13346 "Straight Waveguide" sch_x=55 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6674 N$13347 N$13348 "Straight Waveguide" sch_x=55 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6675 N$13349 N$13350 "Straight Waveguide" sch_x=55 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6676 N$13351 N$13352 "Straight Waveguide" sch_x=55 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6677 N$13353 N$13354 "Straight Waveguide" sch_x=55 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6678 N$13355 N$13356 "Straight Waveguide" sch_x=55 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6679 N$13357 N$13358 "Straight Waveguide" sch_x=55 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6680 N$13359 N$13360 "Straight Waveguide" sch_x=55 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6681 N$13361 N$13362 "Straight Waveguide" sch_x=55 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6682 N$13363 N$13364 "Straight Waveguide" sch_x=55 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6683 N$13365 N$13366 "Straight Waveguide" sch_x=55 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6684 N$13367 N$13368 "Straight Waveguide" sch_x=55 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6685 N$13369 N$13370 "Straight Waveguide" sch_x=53 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6686 N$13371 N$13372 "Straight Waveguide" sch_x=53 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6687 N$13373 N$13374 "Straight Waveguide" sch_x=53 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6688 N$13375 N$13376 "Straight Waveguide" sch_x=53 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6689 N$13377 N$13378 "Straight Waveguide" sch_x=53 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6690 N$13379 N$13380 "Straight Waveguide" sch_x=53 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6691 N$13381 N$13382 "Straight Waveguide" sch_x=53 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6692 N$13383 N$13384 "Straight Waveguide" sch_x=53 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6693 N$13385 N$13386 "Straight Waveguide" sch_x=53 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6694 N$13387 N$13388 "Straight Waveguide" sch_x=53 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6695 N$13389 N$13390 "Straight Waveguide" sch_x=53 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6696 N$13391 N$13392 "Straight Waveguide" sch_x=53 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6697 N$13393 N$13394 "Straight Waveguide" sch_x=53 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6698 N$13395 N$13396 "Straight Waveguide" sch_x=53 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6699 N$13397 N$13398 "Straight Waveguide" sch_x=53 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6700 N$13399 N$13400 "Straight Waveguide" sch_x=53 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6701 N$13401 N$13402 "Straight Waveguide" sch_x=53 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6702 N$13403 N$13404 "Straight Waveguide" sch_x=53 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6703 N$13405 N$13406 "Straight Waveguide" sch_x=53 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6704 N$13407 N$13408 "Straight Waveguide" sch_x=53 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6705 N$13409 N$13410 "Straight Waveguide" sch_x=53 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6706 N$13411 N$13412 "Straight Waveguide" sch_x=53 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6707 N$13413 N$13414 "Straight Waveguide" sch_x=51 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6708 N$13415 N$13416 "Straight Waveguide" sch_x=51 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6709 N$13417 N$13418 "Straight Waveguide" sch_x=51 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6710 N$13419 N$13420 "Straight Waveguide" sch_x=51 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6711 N$13421 N$13422 "Straight Waveguide" sch_x=51 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6712 N$13423 N$13424 "Straight Waveguide" sch_x=51 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6713 N$13425 N$13426 "Straight Waveguide" sch_x=51 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6714 N$13427 N$13428 "Straight Waveguide" sch_x=51 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6715 N$13429 N$13430 "Straight Waveguide" sch_x=51 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6716 N$13431 N$13432 "Straight Waveguide" sch_x=51 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6717 N$13433 N$13434 "Straight Waveguide" sch_x=51 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6718 N$13435 N$13436 "Straight Waveguide" sch_x=51 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6719 N$13437 N$13438 "Straight Waveguide" sch_x=51 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6720 N$13439 N$13440 "Straight Waveguide" sch_x=51 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6721 N$13441 N$13442 "Straight Waveguide" sch_x=51 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6722 N$13443 N$13444 "Straight Waveguide" sch_x=51 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6723 N$13445 N$13446 "Straight Waveguide" sch_x=51 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6724 N$13447 N$13448 "Straight Waveguide" sch_x=51 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6725 N$13449 N$13450 "Straight Waveguide" sch_x=51 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6726 N$13451 N$13452 "Straight Waveguide" sch_x=51 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6727 N$13453 N$13454 "Straight Waveguide" sch_x=49 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6728 N$13455 N$13456 "Straight Waveguide" sch_x=49 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6729 N$13457 N$13458 "Straight Waveguide" sch_x=49 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6730 N$13459 N$13460 "Straight Waveguide" sch_x=49 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6731 N$13461 N$13462 "Straight Waveguide" sch_x=49 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6732 N$13463 N$13464 "Straight Waveguide" sch_x=49 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6733 N$13465 N$13466 "Straight Waveguide" sch_x=49 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6734 N$13467 N$13468 "Straight Waveguide" sch_x=49 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6735 N$13469 N$13470 "Straight Waveguide" sch_x=49 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6736 N$13471 N$13472 "Straight Waveguide" sch_x=49 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6737 N$13473 N$13474 "Straight Waveguide" sch_x=49 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6738 N$13475 N$13476 "Straight Waveguide" sch_x=49 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6739 N$13477 N$13478 "Straight Waveguide" sch_x=49 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6740 N$13479 N$13480 "Straight Waveguide" sch_x=49 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6741 N$13481 N$13482 "Straight Waveguide" sch_x=49 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6742 N$13483 N$13484 "Straight Waveguide" sch_x=49 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6743 N$13485 N$13486 "Straight Waveguide" sch_x=49 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6744 N$13487 N$13488 "Straight Waveguide" sch_x=49 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6745 N$13489 N$13490 "Straight Waveguide" sch_x=47 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6746 N$13491 N$13492 "Straight Waveguide" sch_x=47 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6747 N$13493 N$13494 "Straight Waveguide" sch_x=47 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6748 N$13495 N$13496 "Straight Waveguide" sch_x=47 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6749 N$13497 N$13498 "Straight Waveguide" sch_x=47 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6750 N$13499 N$13500 "Straight Waveguide" sch_x=47 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6751 N$13501 N$13502 "Straight Waveguide" sch_x=47 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6752 N$13503 N$13504 "Straight Waveguide" sch_x=47 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6753 N$13505 N$13506 "Straight Waveguide" sch_x=47 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6754 N$13507 N$13508 "Straight Waveguide" sch_x=47 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6755 N$13509 N$13510 "Straight Waveguide" sch_x=47 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6756 N$13511 N$13512 "Straight Waveguide" sch_x=47 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6757 N$13513 N$13514 "Straight Waveguide" sch_x=47 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6758 N$13515 N$13516 "Straight Waveguide" sch_x=47 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6759 N$13517 N$13518 "Straight Waveguide" sch_x=47 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6760 N$13519 N$13520 "Straight Waveguide" sch_x=47 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6761 N$13521 N$13522 "Straight Waveguide" sch_x=45 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6762 N$13523 N$13524 "Straight Waveguide" sch_x=45 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6763 N$13525 N$13526 "Straight Waveguide" sch_x=45 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6764 N$13527 N$13528 "Straight Waveguide" sch_x=45 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6765 N$13529 N$13530 "Straight Waveguide" sch_x=45 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6766 N$13531 N$13532 "Straight Waveguide" sch_x=45 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6767 N$13533 N$13534 "Straight Waveguide" sch_x=45 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6768 N$13535 N$13536 "Straight Waveguide" sch_x=45 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6769 N$13537 N$13538 "Straight Waveguide" sch_x=45 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6770 N$13539 N$13540 "Straight Waveguide" sch_x=45 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6771 N$13541 N$13542 "Straight Waveguide" sch_x=45 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6772 N$13543 N$13544 "Straight Waveguide" sch_x=45 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6773 N$13545 N$13546 "Straight Waveguide" sch_x=45 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6774 N$13547 N$13548 "Straight Waveguide" sch_x=45 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6775 N$13549 N$13550 "Straight Waveguide" sch_x=43 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6776 N$13551 N$13552 "Straight Waveguide" sch_x=43 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6777 N$13553 N$13554 "Straight Waveguide" sch_x=43 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6778 N$13555 N$13556 "Straight Waveguide" sch_x=43 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6779 N$13557 N$13558 "Straight Waveguide" sch_x=43 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6780 N$13559 N$13560 "Straight Waveguide" sch_x=43 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6781 N$13561 N$13562 "Straight Waveguide" sch_x=43 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6782 N$13563 N$13564 "Straight Waveguide" sch_x=43 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6783 N$13565 N$13566 "Straight Waveguide" sch_x=43 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6784 N$13567 N$13568 "Straight Waveguide" sch_x=43 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6785 N$13569 N$13570 "Straight Waveguide" sch_x=43 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6786 N$13571 N$13572 "Straight Waveguide" sch_x=43 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6787 N$13573 N$13574 "Straight Waveguide" sch_x=41 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6788 N$13575 N$13576 "Straight Waveguide" sch_x=41 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6789 N$13577 N$13578 "Straight Waveguide" sch_x=41 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6790 N$13579 N$13580 "Straight Waveguide" sch_x=41 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6791 N$13581 N$13582 "Straight Waveguide" sch_x=41 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6792 N$13583 N$13584 "Straight Waveguide" sch_x=41 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6793 N$13585 N$13586 "Straight Waveguide" sch_x=41 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6794 N$13587 N$13588 "Straight Waveguide" sch_x=41 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6795 N$13589 N$13590 "Straight Waveguide" sch_x=41 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6796 N$13591 N$13592 "Straight Waveguide" sch_x=41 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6797 N$13593 N$13594 "Straight Waveguide" sch_x=39 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6798 N$13595 N$13596 "Straight Waveguide" sch_x=39 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6799 N$13597 N$13598 "Straight Waveguide" sch_x=39 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6800 N$13599 N$13600 "Straight Waveguide" sch_x=39 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6801 N$13601 N$13602 "Straight Waveguide" sch_x=39 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6802 N$13603 N$13604 "Straight Waveguide" sch_x=39 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6803 N$13605 N$13606 "Straight Waveguide" sch_x=39 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6804 N$13607 N$13608 "Straight Waveguide" sch_x=39 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6805 N$13609 N$13610 "Straight Waveguide" sch_x=37 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6806 N$13611 N$13612 "Straight Waveguide" sch_x=37 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6807 N$13613 N$13614 "Straight Waveguide" sch_x=37 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6808 N$13615 N$13616 "Straight Waveguide" sch_x=37 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6809 N$13617 N$13618 "Straight Waveguide" sch_x=37 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6810 N$13619 N$13620 "Straight Waveguide" sch_x=37 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6811 N$13621 N$13622 "Straight Waveguide" sch_x=35 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6812 N$13623 N$13624 "Straight Waveguide" sch_x=35 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6813 N$13625 N$13626 "Straight Waveguide" sch_x=35 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6814 N$13627 N$13628 "Straight Waveguide" sch_x=35 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6815 N$13629 N$13630 "Straight Waveguide" sch_x=33 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6816 N$13631 N$13632 "Straight Waveguide" sch_x=33 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6817 N$13634 N$13633 "Straight Waveguide" sch_x=45 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6818 N$13636 N$13635 "Straight Waveguide" sch_x=44 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6819 N$13638 N$13637 "Straight Waveguide" sch_x=43 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6820 N$13640 N$13639 "Straight Waveguide" sch_x=42 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6821 N$13642 N$13641 "Straight Waveguide" sch_x=41 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6822 N$13644 N$13643 "Straight Waveguide" sch_x=40 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6823 N$13646 N$13645 "Straight Waveguide" sch_x=39 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6824 N$13648 N$13647 "Straight Waveguide" sch_x=38 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6825 N$13650 N$13649 "Straight Waveguide" sch_x=37 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6826 N$13652 N$13651 "Straight Waveguide" sch_x=36 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6827 N$13654 N$13653 "Straight Waveguide" sch_x=35 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6828 N$13656 N$13655 "Straight Waveguide" sch_x=34 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6829 N$13658 N$13657 "Straight Waveguide" sch_x=33 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6830 N$13660 N$13659 "Straight Waveguide" sch_x=32 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6831 N$13662 N$13661 "Straight Waveguide" sch_x=31 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6832 N$13664 N$13663 "Straight Waveguide" sch_x=31 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6833 N$13666 N$13665 "Straight Waveguide" sch_x=32 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6834 N$13668 N$13667 "Straight Waveguide" sch_x=33 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6835 N$13670 N$13669 "Straight Waveguide" sch_x=34 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6836 N$13672 N$13671 "Straight Waveguide" sch_x=35 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6837 N$13674 N$13673 "Straight Waveguide" sch_x=36 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6838 N$13676 N$13675 "Straight Waveguide" sch_x=37 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6839 N$13678 N$13677 "Straight Waveguide" sch_x=38 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6840 N$13680 N$13679 "Straight Waveguide" sch_x=39 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6841 N$13682 N$13681 "Straight Waveguide" sch_x=40 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6842 N$13684 N$13683 "Straight Waveguide" sch_x=41 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6843 N$13686 N$13685 "Straight Waveguide" sch_x=42 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6844 N$13688 N$13687 "Straight Waveguide" sch_x=43 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6845 N$13690 N$13689 "Straight Waveguide" sch_x=44 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6846 N$13692 N$13691 "Straight Waveguide" sch_x=45 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6847 N$13694 N$13693 "Straight Waveguide" sch_x=46 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6848 N$13696 N$13695 "Straight Waveguide" sch_x=46 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6849 N$13698 N$13697 "Straight Waveguide" sch_x=-125 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6850 N$13700 N$13699 "Straight Waveguide" sch_x=-125 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6851 N$13702 N$13701 "Straight Waveguide" sch_x=-125 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6852 N$13704 N$13703 "Straight Waveguide" sch_x=-125 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6853 N$13706 N$13705 "Straight Waveguide" sch_x=-125 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6854 N$13708 N$13707 "Straight Waveguide" sch_x=-125 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6855 N$13710 N$13709 "Straight Waveguide" sch_x=-125 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6856 N$13712 N$13711 "Straight Waveguide" sch_x=-125 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6857 N$13714 N$13713 "Straight Waveguide" sch_x=-125 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6858 N$13716 N$13715 "Straight Waveguide" sch_x=-125 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6859 N$13718 N$13717 "Straight Waveguide" sch_x=-125 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6860 N$13720 N$13719 "Straight Waveguide" sch_x=-125 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6861 N$13722 N$13721 "Straight Waveguide" sch_x=-125 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6862 N$13724 N$13723 "Straight Waveguide" sch_x=-125 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6863 N$13726 N$13725 "Straight Waveguide" sch_x=-125 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6864 N$13728 N$13727 "Straight Waveguide" sch_x=-125 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6865 N$13730 N$13729 "Straight Waveguide" sch_x=-125 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6866 N$13732 N$13731 "Straight Waveguide" sch_x=-125 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6867 N$13734 N$13733 "Straight Waveguide" sch_x=-125 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6868 N$13736 N$13735 "Straight Waveguide" sch_x=-125 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6869 N$13738 N$13737 "Straight Waveguide" sch_x=-125 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6870 N$13740 N$13739 "Straight Waveguide" sch_x=-125 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6871 N$13742 N$13741 "Straight Waveguide" sch_x=-125 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6872 N$13744 N$13743 "Straight Waveguide" sch_x=-125 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6873 N$13746 N$13745 "Straight Waveguide" sch_x=-125 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6874 N$13748 N$13747 "Straight Waveguide" sch_x=-125 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6875 N$13750 N$13749 "Straight Waveguide" sch_x=-125 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6876 N$13752 N$13751 "Straight Waveguide" sch_x=-125 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6877 N$13754 N$13753 "Straight Waveguide" sch_x=-125 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6878 N$13756 N$13755 "Straight Waveguide" sch_x=-125 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6879 N$13758 N$13757 "Straight Waveguide" sch_x=-125 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6880 N$13760 N$13759 "Straight Waveguide" sch_x=-125 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6881 N$13762 N$13761 "Straight Waveguide" sch_x=-125 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6882 N$13764 N$13763 "Straight Waveguide" sch_x=-125 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6883 N$13766 N$13765 "Straight Waveguide" sch_x=-125 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6884 N$13768 N$13767 "Straight Waveguide" sch_x=-125 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6885 N$13770 N$13769 "Straight Waveguide" sch_x=-125 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6886 N$13772 N$13771 "Straight Waveguide" sch_x=-125 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6887 N$13774 N$13773 "Straight Waveguide" sch_x=-125 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6888 N$13776 N$13775 "Straight Waveguide" sch_x=-125 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6889 N$13778 N$13777 "Straight Waveguide" sch_x=-125 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6890 N$13780 N$13779 "Straight Waveguide" sch_x=-125 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6891 N$13782 N$13781 "Straight Waveguide" sch_x=-125 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6892 N$13784 N$13783 "Straight Waveguide" sch_x=-125 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6893 N$13786 N$13785 "Straight Waveguide" sch_x=-125 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6894 N$13788 N$13787 "Straight Waveguide" sch_x=-125 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6895 N$13790 N$13789 "Straight Waveguide" sch_x=-125 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6896 N$13792 N$13791 "Straight Waveguide" sch_x=-125 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6897 N$13794 N$13793 "Straight Waveguide" sch_x=-125 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6898 N$13796 N$13795 "Straight Waveguide" sch_x=-125 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6899 N$13798 N$13797 "Straight Waveguide" sch_x=-125 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6900 N$13800 N$13799 "Straight Waveguide" sch_x=-125 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6901 N$13802 N$13801 "Straight Waveguide" sch_x=-125 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6902 N$13804 N$13803 "Straight Waveguide" sch_x=-125 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6903 N$13806 N$13805 "Straight Waveguide" sch_x=-125 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6904 N$13808 N$13807 "Straight Waveguide" sch_x=-125 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6905 N$13810 N$13809 "Straight Waveguide" sch_x=-125 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6906 N$13812 N$13811 "Straight Waveguide" sch_x=-125 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6907 N$13814 N$13813 "Straight Waveguide" sch_x=-125 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6908 N$13816 N$13815 "Straight Waveguide" sch_x=-125 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6909 N$13818 N$13817 "Straight Waveguide" sch_x=-125 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6910 N$13820 N$13819 "Straight Waveguide" sch_x=-125 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6911 N$13822 N$13821 "Straight Waveguide" sch_x=-123 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6912 N$13824 N$13823 "Straight Waveguide" sch_x=-123 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6913 N$13826 N$13825 "Straight Waveguide" sch_x=-123 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6914 N$13828 N$13827 "Straight Waveguide" sch_x=-123 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6915 N$13830 N$13829 "Straight Waveguide" sch_x=-123 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6916 N$13832 N$13831 "Straight Waveguide" sch_x=-123 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6917 N$13834 N$13833 "Straight Waveguide" sch_x=-123 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6918 N$13836 N$13835 "Straight Waveguide" sch_x=-123 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6919 N$13838 N$13837 "Straight Waveguide" sch_x=-123 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6920 N$13840 N$13839 "Straight Waveguide" sch_x=-123 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6921 N$13842 N$13841 "Straight Waveguide" sch_x=-123 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6922 N$13844 N$13843 "Straight Waveguide" sch_x=-123 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6923 N$13846 N$13845 "Straight Waveguide" sch_x=-123 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6924 N$13848 N$13847 "Straight Waveguide" sch_x=-123 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6925 N$13850 N$13849 "Straight Waveguide" sch_x=-123 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6926 N$13852 N$13851 "Straight Waveguide" sch_x=-123 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6927 N$13854 N$13853 "Straight Waveguide" sch_x=-123 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6928 N$13856 N$13855 "Straight Waveguide" sch_x=-123 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6929 N$13858 N$13857 "Straight Waveguide" sch_x=-123 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6930 N$13860 N$13859 "Straight Waveguide" sch_x=-123 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6931 N$13862 N$13861 "Straight Waveguide" sch_x=-123 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6932 N$13864 N$13863 "Straight Waveguide" sch_x=-123 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6933 N$13866 N$13865 "Straight Waveguide" sch_x=-123 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6934 N$13868 N$13867 "Straight Waveguide" sch_x=-123 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6935 N$13870 N$13869 "Straight Waveguide" sch_x=-123 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6936 N$13872 N$13871 "Straight Waveguide" sch_x=-123 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6937 N$13874 N$13873 "Straight Waveguide" sch_x=-123 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6938 N$13876 N$13875 "Straight Waveguide" sch_x=-123 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6939 N$13878 N$13877 "Straight Waveguide" sch_x=-123 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6940 N$13880 N$13879 "Straight Waveguide" sch_x=-123 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6941 N$13882 N$13881 "Straight Waveguide" sch_x=-123 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6942 N$13884 N$13883 "Straight Waveguide" sch_x=-123 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6943 N$13886 N$13885 "Straight Waveguide" sch_x=-123 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6944 N$13888 N$13887 "Straight Waveguide" sch_x=-123 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6945 N$13890 N$13889 "Straight Waveguide" sch_x=-123 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6946 N$13892 N$13891 "Straight Waveguide" sch_x=-123 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6947 N$13894 N$13893 "Straight Waveguide" sch_x=-123 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6948 N$13896 N$13895 "Straight Waveguide" sch_x=-123 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6949 N$13898 N$13897 "Straight Waveguide" sch_x=-123 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6950 N$13900 N$13899 "Straight Waveguide" sch_x=-123 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6951 N$13902 N$13901 "Straight Waveguide" sch_x=-123 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6952 N$13904 N$13903 "Straight Waveguide" sch_x=-123 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6953 N$13906 N$13905 "Straight Waveguide" sch_x=-123 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6954 N$13908 N$13907 "Straight Waveguide" sch_x=-123 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6955 N$13910 N$13909 "Straight Waveguide" sch_x=-123 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6956 N$13912 N$13911 "Straight Waveguide" sch_x=-123 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6957 N$13914 N$13913 "Straight Waveguide" sch_x=-123 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6958 N$13916 N$13915 "Straight Waveguide" sch_x=-123 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6959 N$13918 N$13917 "Straight Waveguide" sch_x=-123 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6960 N$13920 N$13919 "Straight Waveguide" sch_x=-123 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6961 N$13922 N$13921 "Straight Waveguide" sch_x=-123 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6962 N$13924 N$13923 "Straight Waveguide" sch_x=-123 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6963 N$13926 N$13925 "Straight Waveguide" sch_x=-123 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6964 N$13928 N$13927 "Straight Waveguide" sch_x=-123 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6965 N$13930 N$13929 "Straight Waveguide" sch_x=-123 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6966 N$13932 N$13931 "Straight Waveguide" sch_x=-123 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6967 N$13934 N$13933 "Straight Waveguide" sch_x=-123 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6968 N$13936 N$13935 "Straight Waveguide" sch_x=-123 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6969 N$13938 N$13937 "Straight Waveguide" sch_x=-123 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6970 N$13940 N$13939 "Straight Waveguide" sch_x=-123 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6971 N$13942 N$13941 "Straight Waveguide" sch_x=-121 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6972 N$13944 N$13943 "Straight Waveguide" sch_x=-121 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6973 N$13946 N$13945 "Straight Waveguide" sch_x=-121 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6974 N$13948 N$13947 "Straight Waveguide" sch_x=-121 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6975 N$13950 N$13949 "Straight Waveguide" sch_x=-121 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6976 N$13952 N$13951 "Straight Waveguide" sch_x=-121 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6977 N$13954 N$13953 "Straight Waveguide" sch_x=-121 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6978 N$13956 N$13955 "Straight Waveguide" sch_x=-121 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6979 N$13958 N$13957 "Straight Waveguide" sch_x=-121 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6980 N$13960 N$13959 "Straight Waveguide" sch_x=-121 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6981 N$13962 N$13961 "Straight Waveguide" sch_x=-121 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6982 N$13964 N$13963 "Straight Waveguide" sch_x=-121 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6983 N$13966 N$13965 "Straight Waveguide" sch_x=-121 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6984 N$13968 N$13967 "Straight Waveguide" sch_x=-121 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6985 N$13970 N$13969 "Straight Waveguide" sch_x=-121 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6986 N$13972 N$13971 "Straight Waveguide" sch_x=-121 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6987 N$13974 N$13973 "Straight Waveguide" sch_x=-121 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6988 N$13976 N$13975 "Straight Waveguide" sch_x=-121 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6989 N$13978 N$13977 "Straight Waveguide" sch_x=-121 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6990 N$13980 N$13979 "Straight Waveguide" sch_x=-121 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6991 N$13982 N$13981 "Straight Waveguide" sch_x=-121 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6992 N$13984 N$13983 "Straight Waveguide" sch_x=-121 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6993 N$13986 N$13985 "Straight Waveguide" sch_x=-121 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6994 N$13988 N$13987 "Straight Waveguide" sch_x=-121 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6995 N$13990 N$13989 "Straight Waveguide" sch_x=-121 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6996 N$13992 N$13991 "Straight Waveguide" sch_x=-121 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6997 N$13994 N$13993 "Straight Waveguide" sch_x=-121 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6998 N$13996 N$13995 "Straight Waveguide" sch_x=-121 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6999 N$13998 N$13997 "Straight Waveguide" sch_x=-121 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7000 N$14000 N$13999 "Straight Waveguide" sch_x=-121 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7001 N$14002 N$14001 "Straight Waveguide" sch_x=-121 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7002 N$14004 N$14003 "Straight Waveguide" sch_x=-121 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7003 N$14006 N$14005 "Straight Waveguide" sch_x=-121 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7004 N$14008 N$14007 "Straight Waveguide" sch_x=-121 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7005 N$14010 N$14009 "Straight Waveguide" sch_x=-121 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7006 N$14012 N$14011 "Straight Waveguide" sch_x=-121 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7007 N$14014 N$14013 "Straight Waveguide" sch_x=-121 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7008 N$14016 N$14015 "Straight Waveguide" sch_x=-121 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7009 N$14018 N$14017 "Straight Waveguide" sch_x=-121 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7010 N$14020 N$14019 "Straight Waveguide" sch_x=-121 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7011 N$14022 N$14021 "Straight Waveguide" sch_x=-121 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7012 N$14024 N$14023 "Straight Waveguide" sch_x=-121 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7013 N$14026 N$14025 "Straight Waveguide" sch_x=-121 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7014 N$14028 N$14027 "Straight Waveguide" sch_x=-121 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7015 N$14030 N$14029 "Straight Waveguide" sch_x=-121 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7016 N$14032 N$14031 "Straight Waveguide" sch_x=-121 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7017 N$14034 N$14033 "Straight Waveguide" sch_x=-121 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7018 N$14036 N$14035 "Straight Waveguide" sch_x=-121 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7019 N$14038 N$14037 "Straight Waveguide" sch_x=-121 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7020 N$14040 N$14039 "Straight Waveguide" sch_x=-121 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7021 N$14042 N$14041 "Straight Waveguide" sch_x=-121 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7022 N$14044 N$14043 "Straight Waveguide" sch_x=-121 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7023 N$14046 N$14045 "Straight Waveguide" sch_x=-121 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7024 N$14048 N$14047 "Straight Waveguide" sch_x=-121 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7025 N$14050 N$14049 "Straight Waveguide" sch_x=-121 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7026 N$14052 N$14051 "Straight Waveguide" sch_x=-121 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7027 N$14054 N$14053 "Straight Waveguide" sch_x=-121 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7028 N$14056 N$14055 "Straight Waveguide" sch_x=-121 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7029 N$14058 N$14057 "Straight Waveguide" sch_x=-119 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7030 N$14060 N$14059 "Straight Waveguide" sch_x=-119 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7031 N$14062 N$14061 "Straight Waveguide" sch_x=-119 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7032 N$14064 N$14063 "Straight Waveguide" sch_x=-119 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7033 N$14066 N$14065 "Straight Waveguide" sch_x=-119 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7034 N$14068 N$14067 "Straight Waveguide" sch_x=-119 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7035 N$14070 N$14069 "Straight Waveguide" sch_x=-119 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7036 N$14072 N$14071 "Straight Waveguide" sch_x=-119 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7037 N$14074 N$14073 "Straight Waveguide" sch_x=-119 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7038 N$14076 N$14075 "Straight Waveguide" sch_x=-119 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7039 N$14078 N$14077 "Straight Waveguide" sch_x=-119 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7040 N$14080 N$14079 "Straight Waveguide" sch_x=-119 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7041 N$14082 N$14081 "Straight Waveguide" sch_x=-119 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7042 N$14084 N$14083 "Straight Waveguide" sch_x=-119 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7043 N$14086 N$14085 "Straight Waveguide" sch_x=-119 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7044 N$14088 N$14087 "Straight Waveguide" sch_x=-119 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7045 N$14090 N$14089 "Straight Waveguide" sch_x=-119 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7046 N$14092 N$14091 "Straight Waveguide" sch_x=-119 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7047 N$14094 N$14093 "Straight Waveguide" sch_x=-119 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7048 N$14096 N$14095 "Straight Waveguide" sch_x=-119 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7049 N$14098 N$14097 "Straight Waveguide" sch_x=-119 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7050 N$14100 N$14099 "Straight Waveguide" sch_x=-119 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7051 N$14102 N$14101 "Straight Waveguide" sch_x=-119 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7052 N$14104 N$14103 "Straight Waveguide" sch_x=-119 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7053 N$14106 N$14105 "Straight Waveguide" sch_x=-119 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7054 N$14108 N$14107 "Straight Waveguide" sch_x=-119 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7055 N$14110 N$14109 "Straight Waveguide" sch_x=-119 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7056 N$14112 N$14111 "Straight Waveguide" sch_x=-119 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7057 N$14114 N$14113 "Straight Waveguide" sch_x=-119 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7058 N$14116 N$14115 "Straight Waveguide" sch_x=-119 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7059 N$14118 N$14117 "Straight Waveguide" sch_x=-119 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7060 N$14120 N$14119 "Straight Waveguide" sch_x=-119 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7061 N$14122 N$14121 "Straight Waveguide" sch_x=-119 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7062 N$14124 N$14123 "Straight Waveguide" sch_x=-119 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7063 N$14126 N$14125 "Straight Waveguide" sch_x=-119 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7064 N$14128 N$14127 "Straight Waveguide" sch_x=-119 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7065 N$14130 N$14129 "Straight Waveguide" sch_x=-119 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7066 N$14132 N$14131 "Straight Waveguide" sch_x=-119 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7067 N$14134 N$14133 "Straight Waveguide" sch_x=-119 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7068 N$14136 N$14135 "Straight Waveguide" sch_x=-119 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7069 N$14138 N$14137 "Straight Waveguide" sch_x=-119 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7070 N$14140 N$14139 "Straight Waveguide" sch_x=-119 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7071 N$14142 N$14141 "Straight Waveguide" sch_x=-119 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7072 N$14144 N$14143 "Straight Waveguide" sch_x=-119 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7073 N$14146 N$14145 "Straight Waveguide" sch_x=-119 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7074 N$14148 N$14147 "Straight Waveguide" sch_x=-119 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7075 N$14150 N$14149 "Straight Waveguide" sch_x=-119 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7076 N$14152 N$14151 "Straight Waveguide" sch_x=-119 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7077 N$14154 N$14153 "Straight Waveguide" sch_x=-119 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7078 N$14156 N$14155 "Straight Waveguide" sch_x=-119 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7079 N$14158 N$14157 "Straight Waveguide" sch_x=-119 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7080 N$14160 N$14159 "Straight Waveguide" sch_x=-119 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7081 N$14162 N$14161 "Straight Waveguide" sch_x=-119 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7082 N$14164 N$14163 "Straight Waveguide" sch_x=-119 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7083 N$14166 N$14165 "Straight Waveguide" sch_x=-119 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7084 N$14168 N$14167 "Straight Waveguide" sch_x=-119 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7085 N$14170 N$14169 "Straight Waveguide" sch_x=-117 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7086 N$14172 N$14171 "Straight Waveguide" sch_x=-117 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7087 N$14174 N$14173 "Straight Waveguide" sch_x=-117 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7088 N$14176 N$14175 "Straight Waveguide" sch_x=-117 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7089 N$14178 N$14177 "Straight Waveguide" sch_x=-117 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7090 N$14180 N$14179 "Straight Waveguide" sch_x=-117 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7091 N$14182 N$14181 "Straight Waveguide" sch_x=-117 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7092 N$14184 N$14183 "Straight Waveguide" sch_x=-117 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7093 N$14186 N$14185 "Straight Waveguide" sch_x=-117 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7094 N$14188 N$14187 "Straight Waveguide" sch_x=-117 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7095 N$14190 N$14189 "Straight Waveguide" sch_x=-117 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7096 N$14192 N$14191 "Straight Waveguide" sch_x=-117 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7097 N$14194 N$14193 "Straight Waveguide" sch_x=-117 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7098 N$14196 N$14195 "Straight Waveguide" sch_x=-117 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7099 N$14198 N$14197 "Straight Waveguide" sch_x=-117 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7100 N$14200 N$14199 "Straight Waveguide" sch_x=-117 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7101 N$14202 N$14201 "Straight Waveguide" sch_x=-117 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7102 N$14204 N$14203 "Straight Waveguide" sch_x=-117 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7103 N$14206 N$14205 "Straight Waveguide" sch_x=-117 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7104 N$14208 N$14207 "Straight Waveguide" sch_x=-117 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7105 N$14210 N$14209 "Straight Waveguide" sch_x=-117 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7106 N$14212 N$14211 "Straight Waveguide" sch_x=-117 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7107 N$14214 N$14213 "Straight Waveguide" sch_x=-117 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7108 N$14216 N$14215 "Straight Waveguide" sch_x=-117 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7109 N$14218 N$14217 "Straight Waveguide" sch_x=-117 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7110 N$14220 N$14219 "Straight Waveguide" sch_x=-117 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7111 N$14222 N$14221 "Straight Waveguide" sch_x=-117 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7112 N$14224 N$14223 "Straight Waveguide" sch_x=-117 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7113 N$14226 N$14225 "Straight Waveguide" sch_x=-117 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7114 N$14228 N$14227 "Straight Waveguide" sch_x=-117 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7115 N$14230 N$14229 "Straight Waveguide" sch_x=-117 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7116 N$14232 N$14231 "Straight Waveguide" sch_x=-117 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7117 N$14234 N$14233 "Straight Waveguide" sch_x=-117 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7118 N$14236 N$14235 "Straight Waveguide" sch_x=-117 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7119 N$14238 N$14237 "Straight Waveguide" sch_x=-117 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7120 N$14240 N$14239 "Straight Waveguide" sch_x=-117 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7121 N$14242 N$14241 "Straight Waveguide" sch_x=-117 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7122 N$14244 N$14243 "Straight Waveguide" sch_x=-117 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7123 N$14246 N$14245 "Straight Waveguide" sch_x=-117 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7124 N$14248 N$14247 "Straight Waveguide" sch_x=-117 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7125 N$14250 N$14249 "Straight Waveguide" sch_x=-117 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7126 N$14252 N$14251 "Straight Waveguide" sch_x=-117 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7127 N$14254 N$14253 "Straight Waveguide" sch_x=-117 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7128 N$14256 N$14255 "Straight Waveguide" sch_x=-117 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7129 N$14258 N$14257 "Straight Waveguide" sch_x=-117 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7130 N$14260 N$14259 "Straight Waveguide" sch_x=-117 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7131 N$14262 N$14261 "Straight Waveguide" sch_x=-117 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7132 N$14264 N$14263 "Straight Waveguide" sch_x=-117 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7133 N$14266 N$14265 "Straight Waveguide" sch_x=-117 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7134 N$14268 N$14267 "Straight Waveguide" sch_x=-117 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7135 N$14270 N$14269 "Straight Waveguide" sch_x=-117 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7136 N$14272 N$14271 "Straight Waveguide" sch_x=-117 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7137 N$14274 N$14273 "Straight Waveguide" sch_x=-117 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7138 N$14276 N$14275 "Straight Waveguide" sch_x=-117 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7139 N$14278 N$14277 "Straight Waveguide" sch_x=-115 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7140 N$14280 N$14279 "Straight Waveguide" sch_x=-115 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7141 N$14282 N$14281 "Straight Waveguide" sch_x=-115 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7142 N$14284 N$14283 "Straight Waveguide" sch_x=-115 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7143 N$14286 N$14285 "Straight Waveguide" sch_x=-115 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7144 N$14288 N$14287 "Straight Waveguide" sch_x=-115 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7145 N$14290 N$14289 "Straight Waveguide" sch_x=-115 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7146 N$14292 N$14291 "Straight Waveguide" sch_x=-115 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7147 N$14294 N$14293 "Straight Waveguide" sch_x=-115 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7148 N$14296 N$14295 "Straight Waveguide" sch_x=-115 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7149 N$14298 N$14297 "Straight Waveguide" sch_x=-115 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7150 N$14300 N$14299 "Straight Waveguide" sch_x=-115 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7151 N$14302 N$14301 "Straight Waveguide" sch_x=-115 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7152 N$14304 N$14303 "Straight Waveguide" sch_x=-115 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7153 N$14306 N$14305 "Straight Waveguide" sch_x=-115 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7154 N$14308 N$14307 "Straight Waveguide" sch_x=-115 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7155 N$14310 N$14309 "Straight Waveguide" sch_x=-115 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7156 N$14312 N$14311 "Straight Waveguide" sch_x=-115 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7157 N$14314 N$14313 "Straight Waveguide" sch_x=-115 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7158 N$14316 N$14315 "Straight Waveguide" sch_x=-115 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7159 N$14318 N$14317 "Straight Waveguide" sch_x=-115 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7160 N$14320 N$14319 "Straight Waveguide" sch_x=-115 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7161 N$14322 N$14321 "Straight Waveguide" sch_x=-115 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7162 N$14324 N$14323 "Straight Waveguide" sch_x=-115 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7163 N$14326 N$14325 "Straight Waveguide" sch_x=-115 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7164 N$14328 N$14327 "Straight Waveguide" sch_x=-115 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7165 N$14330 N$14329 "Straight Waveguide" sch_x=-115 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7166 N$14332 N$14331 "Straight Waveguide" sch_x=-115 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7167 N$14334 N$14333 "Straight Waveguide" sch_x=-115 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7168 N$14336 N$14335 "Straight Waveguide" sch_x=-115 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7169 N$14338 N$14337 "Straight Waveguide" sch_x=-115 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7170 N$14340 N$14339 "Straight Waveguide" sch_x=-115 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7171 N$14342 N$14341 "Straight Waveguide" sch_x=-115 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7172 N$14344 N$14343 "Straight Waveguide" sch_x=-115 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7173 N$14346 N$14345 "Straight Waveguide" sch_x=-115 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7174 N$14348 N$14347 "Straight Waveguide" sch_x=-115 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7175 N$14350 N$14349 "Straight Waveguide" sch_x=-115 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7176 N$14352 N$14351 "Straight Waveguide" sch_x=-115 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7177 N$14354 N$14353 "Straight Waveguide" sch_x=-115 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7178 N$14356 N$14355 "Straight Waveguide" sch_x=-115 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7179 N$14358 N$14357 "Straight Waveguide" sch_x=-115 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7180 N$14360 N$14359 "Straight Waveguide" sch_x=-115 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7181 N$14362 N$14361 "Straight Waveguide" sch_x=-115 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7182 N$14364 N$14363 "Straight Waveguide" sch_x=-115 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7183 N$14366 N$14365 "Straight Waveguide" sch_x=-115 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7184 N$14368 N$14367 "Straight Waveguide" sch_x=-115 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7185 N$14370 N$14369 "Straight Waveguide" sch_x=-115 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7186 N$14372 N$14371 "Straight Waveguide" sch_x=-115 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7187 N$14374 N$14373 "Straight Waveguide" sch_x=-115 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7188 N$14376 N$14375 "Straight Waveguide" sch_x=-115 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7189 N$14378 N$14377 "Straight Waveguide" sch_x=-115 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7190 N$14380 N$14379 "Straight Waveguide" sch_x=-115 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7191 N$14382 N$14381 "Straight Waveguide" sch_x=-113 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7192 N$14384 N$14383 "Straight Waveguide" sch_x=-113 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7193 N$14386 N$14385 "Straight Waveguide" sch_x=-113 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7194 N$14388 N$14387 "Straight Waveguide" sch_x=-113 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7195 N$14390 N$14389 "Straight Waveguide" sch_x=-113 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7196 N$14392 N$14391 "Straight Waveguide" sch_x=-113 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7197 N$14394 N$14393 "Straight Waveguide" sch_x=-113 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7198 N$14396 N$14395 "Straight Waveguide" sch_x=-113 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7199 N$14398 N$14397 "Straight Waveguide" sch_x=-113 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7200 N$14400 N$14399 "Straight Waveguide" sch_x=-113 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7201 N$14402 N$14401 "Straight Waveguide" sch_x=-113 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7202 N$14404 N$14403 "Straight Waveguide" sch_x=-113 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7203 N$14406 N$14405 "Straight Waveguide" sch_x=-113 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7204 N$14408 N$14407 "Straight Waveguide" sch_x=-113 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7205 N$14410 N$14409 "Straight Waveguide" sch_x=-113 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7206 N$14412 N$14411 "Straight Waveguide" sch_x=-113 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7207 N$14414 N$14413 "Straight Waveguide" sch_x=-113 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7208 N$14416 N$14415 "Straight Waveguide" sch_x=-113 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7209 N$14418 N$14417 "Straight Waveguide" sch_x=-113 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7210 N$14420 N$14419 "Straight Waveguide" sch_x=-113 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7211 N$14422 N$14421 "Straight Waveguide" sch_x=-113 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7212 N$14424 N$14423 "Straight Waveguide" sch_x=-113 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7213 N$14426 N$14425 "Straight Waveguide" sch_x=-113 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7214 N$14428 N$14427 "Straight Waveguide" sch_x=-113 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7215 N$14430 N$14429 "Straight Waveguide" sch_x=-113 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7216 N$14432 N$14431 "Straight Waveguide" sch_x=-113 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7217 N$14434 N$14433 "Straight Waveguide" sch_x=-113 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7218 N$14436 N$14435 "Straight Waveguide" sch_x=-113 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7219 N$14438 N$14437 "Straight Waveguide" sch_x=-113 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7220 N$14440 N$14439 "Straight Waveguide" sch_x=-113 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7221 N$14442 N$14441 "Straight Waveguide" sch_x=-113 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7222 N$14444 N$14443 "Straight Waveguide" sch_x=-113 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7223 N$14446 N$14445 "Straight Waveguide" sch_x=-113 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7224 N$14448 N$14447 "Straight Waveguide" sch_x=-113 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7225 N$14450 N$14449 "Straight Waveguide" sch_x=-113 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7226 N$14452 N$14451 "Straight Waveguide" sch_x=-113 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7227 N$14454 N$14453 "Straight Waveguide" sch_x=-113 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7228 N$14456 N$14455 "Straight Waveguide" sch_x=-113 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7229 N$14458 N$14457 "Straight Waveguide" sch_x=-113 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7230 N$14460 N$14459 "Straight Waveguide" sch_x=-113 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7231 N$14462 N$14461 "Straight Waveguide" sch_x=-113 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7232 N$14464 N$14463 "Straight Waveguide" sch_x=-113 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7233 N$14466 N$14465 "Straight Waveguide" sch_x=-113 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7234 N$14468 N$14467 "Straight Waveguide" sch_x=-113 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7235 N$14470 N$14469 "Straight Waveguide" sch_x=-113 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7236 N$14472 N$14471 "Straight Waveguide" sch_x=-113 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7237 N$14474 N$14473 "Straight Waveguide" sch_x=-113 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7238 N$14476 N$14475 "Straight Waveguide" sch_x=-113 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7239 N$14478 N$14477 "Straight Waveguide" sch_x=-113 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7240 N$14480 N$14479 "Straight Waveguide" sch_x=-113 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7241 N$14482 N$14481 "Straight Waveguide" sch_x=-111 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7242 N$14484 N$14483 "Straight Waveguide" sch_x=-111 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7243 N$14486 N$14485 "Straight Waveguide" sch_x=-111 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7244 N$14488 N$14487 "Straight Waveguide" sch_x=-111 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7245 N$14490 N$14489 "Straight Waveguide" sch_x=-111 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7246 N$14492 N$14491 "Straight Waveguide" sch_x=-111 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7247 N$14494 N$14493 "Straight Waveguide" sch_x=-111 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7248 N$14496 N$14495 "Straight Waveguide" sch_x=-111 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7249 N$14498 N$14497 "Straight Waveguide" sch_x=-111 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7250 N$14500 N$14499 "Straight Waveguide" sch_x=-111 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7251 N$14502 N$14501 "Straight Waveguide" sch_x=-111 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7252 N$14504 N$14503 "Straight Waveguide" sch_x=-111 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7253 N$14506 N$14505 "Straight Waveguide" sch_x=-111 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7254 N$14508 N$14507 "Straight Waveguide" sch_x=-111 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7255 N$14510 N$14509 "Straight Waveguide" sch_x=-111 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7256 N$14512 N$14511 "Straight Waveguide" sch_x=-111 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7257 N$14514 N$14513 "Straight Waveguide" sch_x=-111 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7258 N$14516 N$14515 "Straight Waveguide" sch_x=-111 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7259 N$14518 N$14517 "Straight Waveguide" sch_x=-111 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7260 N$14520 N$14519 "Straight Waveguide" sch_x=-111 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7261 N$14522 N$14521 "Straight Waveguide" sch_x=-111 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7262 N$14524 N$14523 "Straight Waveguide" sch_x=-111 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7263 N$14526 N$14525 "Straight Waveguide" sch_x=-111 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7264 N$14528 N$14527 "Straight Waveguide" sch_x=-111 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7265 N$14530 N$14529 "Straight Waveguide" sch_x=-111 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7266 N$14532 N$14531 "Straight Waveguide" sch_x=-111 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7267 N$14534 N$14533 "Straight Waveguide" sch_x=-111 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7268 N$14536 N$14535 "Straight Waveguide" sch_x=-111 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7269 N$14538 N$14537 "Straight Waveguide" sch_x=-111 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7270 N$14540 N$14539 "Straight Waveguide" sch_x=-111 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7271 N$14542 N$14541 "Straight Waveguide" sch_x=-111 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7272 N$14544 N$14543 "Straight Waveguide" sch_x=-111 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7273 N$14546 N$14545 "Straight Waveguide" sch_x=-111 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7274 N$14548 N$14547 "Straight Waveguide" sch_x=-111 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7275 N$14550 N$14549 "Straight Waveguide" sch_x=-111 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7276 N$14552 N$14551 "Straight Waveguide" sch_x=-111 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7277 N$14554 N$14553 "Straight Waveguide" sch_x=-111 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7278 N$14556 N$14555 "Straight Waveguide" sch_x=-111 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7279 N$14558 N$14557 "Straight Waveguide" sch_x=-111 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7280 N$14560 N$14559 "Straight Waveguide" sch_x=-111 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7281 N$14562 N$14561 "Straight Waveguide" sch_x=-111 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7282 N$14564 N$14563 "Straight Waveguide" sch_x=-111 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7283 N$14566 N$14565 "Straight Waveguide" sch_x=-111 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7284 N$14568 N$14567 "Straight Waveguide" sch_x=-111 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7285 N$14570 N$14569 "Straight Waveguide" sch_x=-111 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7286 N$14572 N$14571 "Straight Waveguide" sch_x=-111 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7287 N$14574 N$14573 "Straight Waveguide" sch_x=-111 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7288 N$14576 N$14575 "Straight Waveguide" sch_x=-111 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7289 N$14578 N$14577 "Straight Waveguide" sch_x=-109 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7290 N$14580 N$14579 "Straight Waveguide" sch_x=-109 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7291 N$14582 N$14581 "Straight Waveguide" sch_x=-109 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7292 N$14584 N$14583 "Straight Waveguide" sch_x=-109 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7293 N$14586 N$14585 "Straight Waveguide" sch_x=-109 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7294 N$14588 N$14587 "Straight Waveguide" sch_x=-109 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7295 N$14590 N$14589 "Straight Waveguide" sch_x=-109 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7296 N$14592 N$14591 "Straight Waveguide" sch_x=-109 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7297 N$14594 N$14593 "Straight Waveguide" sch_x=-109 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7298 N$14596 N$14595 "Straight Waveguide" sch_x=-109 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7299 N$14598 N$14597 "Straight Waveguide" sch_x=-109 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7300 N$14600 N$14599 "Straight Waveguide" sch_x=-109 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7301 N$14602 N$14601 "Straight Waveguide" sch_x=-109 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7302 N$14604 N$14603 "Straight Waveguide" sch_x=-109 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7303 N$14606 N$14605 "Straight Waveguide" sch_x=-109 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7304 N$14608 N$14607 "Straight Waveguide" sch_x=-109 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7305 N$14610 N$14609 "Straight Waveguide" sch_x=-109 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7306 N$14612 N$14611 "Straight Waveguide" sch_x=-109 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7307 N$14614 N$14613 "Straight Waveguide" sch_x=-109 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7308 N$14616 N$14615 "Straight Waveguide" sch_x=-109 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7309 N$14618 N$14617 "Straight Waveguide" sch_x=-109 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7310 N$14620 N$14619 "Straight Waveguide" sch_x=-109 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7311 N$14622 N$14621 "Straight Waveguide" sch_x=-109 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7312 N$14624 N$14623 "Straight Waveguide" sch_x=-109 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7313 N$14626 N$14625 "Straight Waveguide" sch_x=-109 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7314 N$14628 N$14627 "Straight Waveguide" sch_x=-109 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7315 N$14630 N$14629 "Straight Waveguide" sch_x=-109 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7316 N$14632 N$14631 "Straight Waveguide" sch_x=-109 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7317 N$14634 N$14633 "Straight Waveguide" sch_x=-109 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7318 N$14636 N$14635 "Straight Waveguide" sch_x=-109 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7319 N$14638 N$14637 "Straight Waveguide" sch_x=-109 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7320 N$14640 N$14639 "Straight Waveguide" sch_x=-109 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7321 N$14642 N$14641 "Straight Waveguide" sch_x=-109 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7322 N$14644 N$14643 "Straight Waveguide" sch_x=-109 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7323 N$14646 N$14645 "Straight Waveguide" sch_x=-109 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7324 N$14648 N$14647 "Straight Waveguide" sch_x=-109 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7325 N$14650 N$14649 "Straight Waveguide" sch_x=-109 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7326 N$14652 N$14651 "Straight Waveguide" sch_x=-109 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7327 N$14654 N$14653 "Straight Waveguide" sch_x=-109 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7328 N$14656 N$14655 "Straight Waveguide" sch_x=-109 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7329 N$14658 N$14657 "Straight Waveguide" sch_x=-109 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7330 N$14660 N$14659 "Straight Waveguide" sch_x=-109 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7331 N$14662 N$14661 "Straight Waveguide" sch_x=-109 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7332 N$14664 N$14663 "Straight Waveguide" sch_x=-109 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7333 N$14666 N$14665 "Straight Waveguide" sch_x=-109 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7334 N$14668 N$14667 "Straight Waveguide" sch_x=-109 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7335 N$14670 N$14669 "Straight Waveguide" sch_x=-107 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7336 N$14672 N$14671 "Straight Waveguide" sch_x=-107 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7337 N$14674 N$14673 "Straight Waveguide" sch_x=-107 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7338 N$14676 N$14675 "Straight Waveguide" sch_x=-107 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7339 N$14678 N$14677 "Straight Waveguide" sch_x=-107 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7340 N$14680 N$14679 "Straight Waveguide" sch_x=-107 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7341 N$14682 N$14681 "Straight Waveguide" sch_x=-107 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7342 N$14684 N$14683 "Straight Waveguide" sch_x=-107 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7343 N$14686 N$14685 "Straight Waveguide" sch_x=-107 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7344 N$14688 N$14687 "Straight Waveguide" sch_x=-107 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7345 N$14690 N$14689 "Straight Waveguide" sch_x=-107 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7346 N$14692 N$14691 "Straight Waveguide" sch_x=-107 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7347 N$14694 N$14693 "Straight Waveguide" sch_x=-107 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7348 N$14696 N$14695 "Straight Waveguide" sch_x=-107 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7349 N$14698 N$14697 "Straight Waveguide" sch_x=-107 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7350 N$14700 N$14699 "Straight Waveguide" sch_x=-107 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7351 N$14702 N$14701 "Straight Waveguide" sch_x=-107 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7352 N$14704 N$14703 "Straight Waveguide" sch_x=-107 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7353 N$14706 N$14705 "Straight Waveguide" sch_x=-107 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7354 N$14708 N$14707 "Straight Waveguide" sch_x=-107 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7355 N$14710 N$14709 "Straight Waveguide" sch_x=-107 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7356 N$14712 N$14711 "Straight Waveguide" sch_x=-107 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7357 N$14714 N$14713 "Straight Waveguide" sch_x=-107 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7358 N$14716 N$14715 "Straight Waveguide" sch_x=-107 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7359 N$14718 N$14717 "Straight Waveguide" sch_x=-107 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7360 N$14720 N$14719 "Straight Waveguide" sch_x=-107 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7361 N$14722 N$14721 "Straight Waveguide" sch_x=-107 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7362 N$14724 N$14723 "Straight Waveguide" sch_x=-107 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7363 N$14726 N$14725 "Straight Waveguide" sch_x=-107 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7364 N$14728 N$14727 "Straight Waveguide" sch_x=-107 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7365 N$14730 N$14729 "Straight Waveguide" sch_x=-107 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7366 N$14732 N$14731 "Straight Waveguide" sch_x=-107 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7367 N$14734 N$14733 "Straight Waveguide" sch_x=-107 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7368 N$14736 N$14735 "Straight Waveguide" sch_x=-107 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7369 N$14738 N$14737 "Straight Waveguide" sch_x=-107 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7370 N$14740 N$14739 "Straight Waveguide" sch_x=-107 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7371 N$14742 N$14741 "Straight Waveguide" sch_x=-107 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7372 N$14744 N$14743 "Straight Waveguide" sch_x=-107 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7373 N$14746 N$14745 "Straight Waveguide" sch_x=-107 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7374 N$14748 N$14747 "Straight Waveguide" sch_x=-107 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7375 N$14750 N$14749 "Straight Waveguide" sch_x=-107 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7376 N$14752 N$14751 "Straight Waveguide" sch_x=-107 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7377 N$14754 N$14753 "Straight Waveguide" sch_x=-107 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7378 N$14756 N$14755 "Straight Waveguide" sch_x=-107 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7379 N$14758 N$14757 "Straight Waveguide" sch_x=-105 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7380 N$14760 N$14759 "Straight Waveguide" sch_x=-105 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7381 N$14762 N$14761 "Straight Waveguide" sch_x=-105 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7382 N$14764 N$14763 "Straight Waveguide" sch_x=-105 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7383 N$14766 N$14765 "Straight Waveguide" sch_x=-105 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7384 N$14768 N$14767 "Straight Waveguide" sch_x=-105 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7385 N$14770 N$14769 "Straight Waveguide" sch_x=-105 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7386 N$14772 N$14771 "Straight Waveguide" sch_x=-105 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7387 N$14774 N$14773 "Straight Waveguide" sch_x=-105 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7388 N$14776 N$14775 "Straight Waveguide" sch_x=-105 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7389 N$14778 N$14777 "Straight Waveguide" sch_x=-105 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7390 N$14780 N$14779 "Straight Waveguide" sch_x=-105 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7391 N$14782 N$14781 "Straight Waveguide" sch_x=-105 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7392 N$14784 N$14783 "Straight Waveguide" sch_x=-105 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7393 N$14786 N$14785 "Straight Waveguide" sch_x=-105 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7394 N$14788 N$14787 "Straight Waveguide" sch_x=-105 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7395 N$14790 N$14789 "Straight Waveguide" sch_x=-105 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7396 N$14792 N$14791 "Straight Waveguide" sch_x=-105 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7397 N$14794 N$14793 "Straight Waveguide" sch_x=-105 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7398 N$14796 N$14795 "Straight Waveguide" sch_x=-105 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7399 N$14798 N$14797 "Straight Waveguide" sch_x=-105 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7400 N$14800 N$14799 "Straight Waveguide" sch_x=-105 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7401 N$14802 N$14801 "Straight Waveguide" sch_x=-105 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7402 N$14804 N$14803 "Straight Waveguide" sch_x=-105 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7403 N$14806 N$14805 "Straight Waveguide" sch_x=-105 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7404 N$14808 N$14807 "Straight Waveguide" sch_x=-105 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7405 N$14810 N$14809 "Straight Waveguide" sch_x=-105 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7406 N$14812 N$14811 "Straight Waveguide" sch_x=-105 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7407 N$14814 N$14813 "Straight Waveguide" sch_x=-105 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7408 N$14816 N$14815 "Straight Waveguide" sch_x=-105 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7409 N$14818 N$14817 "Straight Waveguide" sch_x=-105 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7410 N$14820 N$14819 "Straight Waveguide" sch_x=-105 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7411 N$14822 N$14821 "Straight Waveguide" sch_x=-105 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7412 N$14824 N$14823 "Straight Waveguide" sch_x=-105 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7413 N$14826 N$14825 "Straight Waveguide" sch_x=-105 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7414 N$14828 N$14827 "Straight Waveguide" sch_x=-105 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7415 N$14830 N$14829 "Straight Waveguide" sch_x=-105 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7416 N$14832 N$14831 "Straight Waveguide" sch_x=-105 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7417 N$14834 N$14833 "Straight Waveguide" sch_x=-105 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7418 N$14836 N$14835 "Straight Waveguide" sch_x=-105 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7419 N$14838 N$14837 "Straight Waveguide" sch_x=-105 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7420 N$14840 N$14839 "Straight Waveguide" sch_x=-105 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7421 N$14842 N$14841 "Straight Waveguide" sch_x=-103 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7422 N$14844 N$14843 "Straight Waveguide" sch_x=-103 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7423 N$14846 N$14845 "Straight Waveguide" sch_x=-103 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7424 N$14848 N$14847 "Straight Waveguide" sch_x=-103 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7425 N$14850 N$14849 "Straight Waveguide" sch_x=-103 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7426 N$14852 N$14851 "Straight Waveguide" sch_x=-103 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7427 N$14854 N$14853 "Straight Waveguide" sch_x=-103 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7428 N$14856 N$14855 "Straight Waveguide" sch_x=-103 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7429 N$14858 N$14857 "Straight Waveguide" sch_x=-103 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7430 N$14860 N$14859 "Straight Waveguide" sch_x=-103 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7431 N$14862 N$14861 "Straight Waveguide" sch_x=-103 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7432 N$14864 N$14863 "Straight Waveguide" sch_x=-103 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7433 N$14866 N$14865 "Straight Waveguide" sch_x=-103 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7434 N$14868 N$14867 "Straight Waveguide" sch_x=-103 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7435 N$14870 N$14869 "Straight Waveguide" sch_x=-103 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7436 N$14872 N$14871 "Straight Waveguide" sch_x=-103 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7437 N$14874 N$14873 "Straight Waveguide" sch_x=-103 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7438 N$14876 N$14875 "Straight Waveguide" sch_x=-103 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7439 N$14878 N$14877 "Straight Waveguide" sch_x=-103 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7440 N$14880 N$14879 "Straight Waveguide" sch_x=-103 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7441 N$14882 N$14881 "Straight Waveguide" sch_x=-103 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7442 N$14884 N$14883 "Straight Waveguide" sch_x=-103 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7443 N$14886 N$14885 "Straight Waveguide" sch_x=-103 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7444 N$14888 N$14887 "Straight Waveguide" sch_x=-103 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7445 N$14890 N$14889 "Straight Waveguide" sch_x=-103 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7446 N$14892 N$14891 "Straight Waveguide" sch_x=-103 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7447 N$14894 N$14893 "Straight Waveguide" sch_x=-103 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7448 N$14896 N$14895 "Straight Waveguide" sch_x=-103 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7449 N$14898 N$14897 "Straight Waveguide" sch_x=-103 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7450 N$14900 N$14899 "Straight Waveguide" sch_x=-103 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7451 N$14902 N$14901 "Straight Waveguide" sch_x=-103 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7452 N$14904 N$14903 "Straight Waveguide" sch_x=-103 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7453 N$14906 N$14905 "Straight Waveguide" sch_x=-103 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7454 N$14908 N$14907 "Straight Waveguide" sch_x=-103 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7455 N$14910 N$14909 "Straight Waveguide" sch_x=-103 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7456 N$14912 N$14911 "Straight Waveguide" sch_x=-103 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7457 N$14914 N$14913 "Straight Waveguide" sch_x=-103 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7458 N$14916 N$14915 "Straight Waveguide" sch_x=-103 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7459 N$14918 N$14917 "Straight Waveguide" sch_x=-103 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7460 N$14920 N$14919 "Straight Waveguide" sch_x=-103 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7461 N$14922 N$14921 "Straight Waveguide" sch_x=-101 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7462 N$14924 N$14923 "Straight Waveguide" sch_x=-101 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7463 N$14926 N$14925 "Straight Waveguide" sch_x=-101 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7464 N$14928 N$14927 "Straight Waveguide" sch_x=-101 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7465 N$14930 N$14929 "Straight Waveguide" sch_x=-101 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7466 N$14932 N$14931 "Straight Waveguide" sch_x=-101 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7467 N$14934 N$14933 "Straight Waveguide" sch_x=-101 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7468 N$14936 N$14935 "Straight Waveguide" sch_x=-101 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7469 N$14938 N$14937 "Straight Waveguide" sch_x=-101 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7470 N$14940 N$14939 "Straight Waveguide" sch_x=-101 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7471 N$14942 N$14941 "Straight Waveguide" sch_x=-101 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7472 N$14944 N$14943 "Straight Waveguide" sch_x=-101 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7473 N$14946 N$14945 "Straight Waveguide" sch_x=-101 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7474 N$14948 N$14947 "Straight Waveguide" sch_x=-101 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7475 N$14950 N$14949 "Straight Waveguide" sch_x=-101 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7476 N$14952 N$14951 "Straight Waveguide" sch_x=-101 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7477 N$14954 N$14953 "Straight Waveguide" sch_x=-101 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7478 N$14956 N$14955 "Straight Waveguide" sch_x=-101 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7479 N$14958 N$14957 "Straight Waveguide" sch_x=-101 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7480 N$14960 N$14959 "Straight Waveguide" sch_x=-101 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7481 N$14962 N$14961 "Straight Waveguide" sch_x=-101 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7482 N$14964 N$14963 "Straight Waveguide" sch_x=-101 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7483 N$14966 N$14965 "Straight Waveguide" sch_x=-101 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7484 N$14968 N$14967 "Straight Waveguide" sch_x=-101 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7485 N$14970 N$14969 "Straight Waveguide" sch_x=-101 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7486 N$14972 N$14971 "Straight Waveguide" sch_x=-101 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7487 N$14974 N$14973 "Straight Waveguide" sch_x=-101 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7488 N$14976 N$14975 "Straight Waveguide" sch_x=-101 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7489 N$14978 N$14977 "Straight Waveguide" sch_x=-101 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7490 N$14980 N$14979 "Straight Waveguide" sch_x=-101 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7491 N$14982 N$14981 "Straight Waveguide" sch_x=-101 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7492 N$14984 N$14983 "Straight Waveguide" sch_x=-101 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7493 N$14986 N$14985 "Straight Waveguide" sch_x=-101 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7494 N$14988 N$14987 "Straight Waveguide" sch_x=-101 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7495 N$14990 N$14989 "Straight Waveguide" sch_x=-101 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7496 N$14992 N$14991 "Straight Waveguide" sch_x=-101 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7497 N$14994 N$14993 "Straight Waveguide" sch_x=-101 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7498 N$14996 N$14995 "Straight Waveguide" sch_x=-101 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7499 N$14998 N$14997 "Straight Waveguide" sch_x=-99 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7500 N$15000 N$14999 "Straight Waveguide" sch_x=-99 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7501 N$15002 N$15001 "Straight Waveguide" sch_x=-99 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7502 N$15004 N$15003 "Straight Waveguide" sch_x=-99 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7503 N$15006 N$15005 "Straight Waveguide" sch_x=-99 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7504 N$15008 N$15007 "Straight Waveguide" sch_x=-99 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7505 N$15010 N$15009 "Straight Waveguide" sch_x=-99 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7506 N$15012 N$15011 "Straight Waveguide" sch_x=-99 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7507 N$15014 N$15013 "Straight Waveguide" sch_x=-99 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7508 N$15016 N$15015 "Straight Waveguide" sch_x=-99 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7509 N$15018 N$15017 "Straight Waveguide" sch_x=-99 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7510 N$15020 N$15019 "Straight Waveguide" sch_x=-99 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7511 N$15022 N$15021 "Straight Waveguide" sch_x=-99 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7512 N$15024 N$15023 "Straight Waveguide" sch_x=-99 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7513 N$15026 N$15025 "Straight Waveguide" sch_x=-99 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7514 N$15028 N$15027 "Straight Waveguide" sch_x=-99 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7515 N$15030 N$15029 "Straight Waveguide" sch_x=-99 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7516 N$15032 N$15031 "Straight Waveguide" sch_x=-99 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7517 N$15034 N$15033 "Straight Waveguide" sch_x=-99 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7518 N$15036 N$15035 "Straight Waveguide" sch_x=-99 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7519 N$15038 N$15037 "Straight Waveguide" sch_x=-99 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7520 N$15040 N$15039 "Straight Waveguide" sch_x=-99 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7521 N$15042 N$15041 "Straight Waveguide" sch_x=-99 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7522 N$15044 N$15043 "Straight Waveguide" sch_x=-99 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7523 N$15046 N$15045 "Straight Waveguide" sch_x=-99 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7524 N$15048 N$15047 "Straight Waveguide" sch_x=-99 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7525 N$15050 N$15049 "Straight Waveguide" sch_x=-99 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7526 N$15052 N$15051 "Straight Waveguide" sch_x=-99 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7527 N$15054 N$15053 "Straight Waveguide" sch_x=-99 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7528 N$15056 N$15055 "Straight Waveguide" sch_x=-99 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7529 N$15058 N$15057 "Straight Waveguide" sch_x=-99 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7530 N$15060 N$15059 "Straight Waveguide" sch_x=-99 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7531 N$15062 N$15061 "Straight Waveguide" sch_x=-99 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7532 N$15064 N$15063 "Straight Waveguide" sch_x=-99 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7533 N$15066 N$15065 "Straight Waveguide" sch_x=-99 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7534 N$15068 N$15067 "Straight Waveguide" sch_x=-99 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7535 N$15070 N$15069 "Straight Waveguide" sch_x=-97 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7536 N$15072 N$15071 "Straight Waveguide" sch_x=-97 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7537 N$15074 N$15073 "Straight Waveguide" sch_x=-97 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7538 N$15076 N$15075 "Straight Waveguide" sch_x=-97 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7539 N$15078 N$15077 "Straight Waveguide" sch_x=-97 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7540 N$15080 N$15079 "Straight Waveguide" sch_x=-97 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7541 N$15082 N$15081 "Straight Waveguide" sch_x=-97 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7542 N$15084 N$15083 "Straight Waveguide" sch_x=-97 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7543 N$15086 N$15085 "Straight Waveguide" sch_x=-97 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7544 N$15088 N$15087 "Straight Waveguide" sch_x=-97 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7545 N$15090 N$15089 "Straight Waveguide" sch_x=-97 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7546 N$15092 N$15091 "Straight Waveguide" sch_x=-97 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7547 N$15094 N$15093 "Straight Waveguide" sch_x=-97 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7548 N$15096 N$15095 "Straight Waveguide" sch_x=-97 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7549 N$15098 N$15097 "Straight Waveguide" sch_x=-97 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7550 N$15100 N$15099 "Straight Waveguide" sch_x=-97 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7551 N$15102 N$15101 "Straight Waveguide" sch_x=-97 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7552 N$15104 N$15103 "Straight Waveguide" sch_x=-97 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7553 N$15106 N$15105 "Straight Waveguide" sch_x=-97 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7554 N$15108 N$15107 "Straight Waveguide" sch_x=-97 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7555 N$15110 N$15109 "Straight Waveguide" sch_x=-97 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7556 N$15112 N$15111 "Straight Waveguide" sch_x=-97 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7557 N$15114 N$15113 "Straight Waveguide" sch_x=-97 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7558 N$15116 N$15115 "Straight Waveguide" sch_x=-97 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7559 N$15118 N$15117 "Straight Waveguide" sch_x=-97 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7560 N$15120 N$15119 "Straight Waveguide" sch_x=-97 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7561 N$15122 N$15121 "Straight Waveguide" sch_x=-97 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7562 N$15124 N$15123 "Straight Waveguide" sch_x=-97 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7563 N$15126 N$15125 "Straight Waveguide" sch_x=-97 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7564 N$15128 N$15127 "Straight Waveguide" sch_x=-97 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7565 N$15130 N$15129 "Straight Waveguide" sch_x=-97 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7566 N$15132 N$15131 "Straight Waveguide" sch_x=-97 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7567 N$15134 N$15133 "Straight Waveguide" sch_x=-97 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7568 N$15136 N$15135 "Straight Waveguide" sch_x=-97 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7569 N$15138 N$15137 "Straight Waveguide" sch_x=-95 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7570 N$15140 N$15139 "Straight Waveguide" sch_x=-95 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7571 N$15142 N$15141 "Straight Waveguide" sch_x=-95 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7572 N$15144 N$15143 "Straight Waveguide" sch_x=-95 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7573 N$15146 N$15145 "Straight Waveguide" sch_x=-95 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7574 N$15148 N$15147 "Straight Waveguide" sch_x=-95 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7575 N$15150 N$15149 "Straight Waveguide" sch_x=-95 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7576 N$15152 N$15151 "Straight Waveguide" sch_x=-95 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7577 N$15154 N$15153 "Straight Waveguide" sch_x=-95 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7578 N$15156 N$15155 "Straight Waveguide" sch_x=-95 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7579 N$15158 N$15157 "Straight Waveguide" sch_x=-95 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7580 N$15160 N$15159 "Straight Waveguide" sch_x=-95 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7581 N$15162 N$15161 "Straight Waveguide" sch_x=-95 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7582 N$15164 N$15163 "Straight Waveguide" sch_x=-95 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7583 N$15166 N$15165 "Straight Waveguide" sch_x=-95 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7584 N$15168 N$15167 "Straight Waveguide" sch_x=-95 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7585 N$15170 N$15169 "Straight Waveguide" sch_x=-95 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7586 N$15172 N$15171 "Straight Waveguide" sch_x=-95 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7587 N$15174 N$15173 "Straight Waveguide" sch_x=-95 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7588 N$15176 N$15175 "Straight Waveguide" sch_x=-95 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7589 N$15178 N$15177 "Straight Waveguide" sch_x=-95 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7590 N$15180 N$15179 "Straight Waveguide" sch_x=-95 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7591 N$15182 N$15181 "Straight Waveguide" sch_x=-95 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7592 N$15184 N$15183 "Straight Waveguide" sch_x=-95 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7593 N$15186 N$15185 "Straight Waveguide" sch_x=-95 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7594 N$15188 N$15187 "Straight Waveguide" sch_x=-95 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7595 N$15190 N$15189 "Straight Waveguide" sch_x=-95 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7596 N$15192 N$15191 "Straight Waveguide" sch_x=-95 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7597 N$15194 N$15193 "Straight Waveguide" sch_x=-95 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7598 N$15196 N$15195 "Straight Waveguide" sch_x=-95 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7599 N$15198 N$15197 "Straight Waveguide" sch_x=-95 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7600 N$15200 N$15199 "Straight Waveguide" sch_x=-95 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7601 N$15202 N$15201 "Straight Waveguide" sch_x=-93 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7602 N$15204 N$15203 "Straight Waveguide" sch_x=-93 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7603 N$15206 N$15205 "Straight Waveguide" sch_x=-93 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7604 N$15208 N$15207 "Straight Waveguide" sch_x=-93 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7605 N$15210 N$15209 "Straight Waveguide" sch_x=-93 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7606 N$15212 N$15211 "Straight Waveguide" sch_x=-93 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7607 N$15214 N$15213 "Straight Waveguide" sch_x=-93 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7608 N$15216 N$15215 "Straight Waveguide" sch_x=-93 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7609 N$15218 N$15217 "Straight Waveguide" sch_x=-93 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7610 N$15220 N$15219 "Straight Waveguide" sch_x=-93 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7611 N$15222 N$15221 "Straight Waveguide" sch_x=-93 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7612 N$15224 N$15223 "Straight Waveguide" sch_x=-93 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7613 N$15226 N$15225 "Straight Waveguide" sch_x=-93 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7614 N$15228 N$15227 "Straight Waveguide" sch_x=-93 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7615 N$15230 N$15229 "Straight Waveguide" sch_x=-93 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7616 N$15232 N$15231 "Straight Waveguide" sch_x=-93 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7617 N$15234 N$15233 "Straight Waveguide" sch_x=-93 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7618 N$15236 N$15235 "Straight Waveguide" sch_x=-93 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7619 N$15238 N$15237 "Straight Waveguide" sch_x=-93 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7620 N$15240 N$15239 "Straight Waveguide" sch_x=-93 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7621 N$15242 N$15241 "Straight Waveguide" sch_x=-93 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7622 N$15244 N$15243 "Straight Waveguide" sch_x=-93 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7623 N$15246 N$15245 "Straight Waveguide" sch_x=-93 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7624 N$15248 N$15247 "Straight Waveguide" sch_x=-93 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7625 N$15250 N$15249 "Straight Waveguide" sch_x=-93 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7626 N$15252 N$15251 "Straight Waveguide" sch_x=-93 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7627 N$15254 N$15253 "Straight Waveguide" sch_x=-93 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7628 N$15256 N$15255 "Straight Waveguide" sch_x=-93 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7629 N$15258 N$15257 "Straight Waveguide" sch_x=-93 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7630 N$15260 N$15259 "Straight Waveguide" sch_x=-93 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7631 N$15262 N$15261 "Straight Waveguide" sch_x=-91 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7632 N$15264 N$15263 "Straight Waveguide" sch_x=-91 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7633 N$15266 N$15265 "Straight Waveguide" sch_x=-91 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7634 N$15268 N$15267 "Straight Waveguide" sch_x=-91 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7635 N$15270 N$15269 "Straight Waveguide" sch_x=-91 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7636 N$15272 N$15271 "Straight Waveguide" sch_x=-91 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7637 N$15274 N$15273 "Straight Waveguide" sch_x=-91 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7638 N$15276 N$15275 "Straight Waveguide" sch_x=-91 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7639 N$15278 N$15277 "Straight Waveguide" sch_x=-91 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7640 N$15280 N$15279 "Straight Waveguide" sch_x=-91 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7641 N$15282 N$15281 "Straight Waveguide" sch_x=-91 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7642 N$15284 N$15283 "Straight Waveguide" sch_x=-91 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7643 N$15286 N$15285 "Straight Waveguide" sch_x=-91 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7644 N$15288 N$15287 "Straight Waveguide" sch_x=-91 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7645 N$15290 N$15289 "Straight Waveguide" sch_x=-91 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7646 N$15292 N$15291 "Straight Waveguide" sch_x=-91 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7647 N$15294 N$15293 "Straight Waveguide" sch_x=-91 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7648 N$15296 N$15295 "Straight Waveguide" sch_x=-91 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7649 N$15298 N$15297 "Straight Waveguide" sch_x=-91 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7650 N$15300 N$15299 "Straight Waveguide" sch_x=-91 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7651 N$15302 N$15301 "Straight Waveguide" sch_x=-91 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7652 N$15304 N$15303 "Straight Waveguide" sch_x=-91 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7653 N$15306 N$15305 "Straight Waveguide" sch_x=-91 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7654 N$15308 N$15307 "Straight Waveguide" sch_x=-91 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7655 N$15310 N$15309 "Straight Waveguide" sch_x=-91 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7656 N$15312 N$15311 "Straight Waveguide" sch_x=-91 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7657 N$15314 N$15313 "Straight Waveguide" sch_x=-91 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7658 N$15316 N$15315 "Straight Waveguide" sch_x=-91 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7659 N$15318 N$15317 "Straight Waveguide" sch_x=-89 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7660 N$15320 N$15319 "Straight Waveguide" sch_x=-89 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7661 N$15322 N$15321 "Straight Waveguide" sch_x=-89 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7662 N$15324 N$15323 "Straight Waveguide" sch_x=-89 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7663 N$15326 N$15325 "Straight Waveguide" sch_x=-89 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7664 N$15328 N$15327 "Straight Waveguide" sch_x=-89 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7665 N$15330 N$15329 "Straight Waveguide" sch_x=-89 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7666 N$15332 N$15331 "Straight Waveguide" sch_x=-89 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7667 N$15334 N$15333 "Straight Waveguide" sch_x=-89 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7668 N$15336 N$15335 "Straight Waveguide" sch_x=-89 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7669 N$15338 N$15337 "Straight Waveguide" sch_x=-89 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7670 N$15340 N$15339 "Straight Waveguide" sch_x=-89 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7671 N$15342 N$15341 "Straight Waveguide" sch_x=-89 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7672 N$15344 N$15343 "Straight Waveguide" sch_x=-89 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7673 N$15346 N$15345 "Straight Waveguide" sch_x=-89 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7674 N$15348 N$15347 "Straight Waveguide" sch_x=-89 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7675 N$15350 N$15349 "Straight Waveguide" sch_x=-89 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7676 N$15352 N$15351 "Straight Waveguide" sch_x=-89 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7677 N$15354 N$15353 "Straight Waveguide" sch_x=-89 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7678 N$15356 N$15355 "Straight Waveguide" sch_x=-89 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7679 N$15358 N$15357 "Straight Waveguide" sch_x=-89 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7680 N$15360 N$15359 "Straight Waveguide" sch_x=-89 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7681 N$15362 N$15361 "Straight Waveguide" sch_x=-89 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7682 N$15364 N$15363 "Straight Waveguide" sch_x=-89 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7683 N$15366 N$15365 "Straight Waveguide" sch_x=-89 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7684 N$15368 N$15367 "Straight Waveguide" sch_x=-89 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7685 N$15370 N$15369 "Straight Waveguide" sch_x=-87 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7686 N$15372 N$15371 "Straight Waveguide" sch_x=-87 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7687 N$15374 N$15373 "Straight Waveguide" sch_x=-87 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7688 N$15376 N$15375 "Straight Waveguide" sch_x=-87 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7689 N$15378 N$15377 "Straight Waveguide" sch_x=-87 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7690 N$15380 N$15379 "Straight Waveguide" sch_x=-87 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7691 N$15382 N$15381 "Straight Waveguide" sch_x=-87 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7692 N$15384 N$15383 "Straight Waveguide" sch_x=-87 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7693 N$15386 N$15385 "Straight Waveguide" sch_x=-87 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7694 N$15388 N$15387 "Straight Waveguide" sch_x=-87 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7695 N$15390 N$15389 "Straight Waveguide" sch_x=-87 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7696 N$15392 N$15391 "Straight Waveguide" sch_x=-87 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7697 N$15394 N$15393 "Straight Waveguide" sch_x=-87 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7698 N$15396 N$15395 "Straight Waveguide" sch_x=-87 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7699 N$15398 N$15397 "Straight Waveguide" sch_x=-87 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7700 N$15400 N$15399 "Straight Waveguide" sch_x=-87 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7701 N$15402 N$15401 "Straight Waveguide" sch_x=-87 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7702 N$15404 N$15403 "Straight Waveguide" sch_x=-87 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7703 N$15406 N$15405 "Straight Waveguide" sch_x=-87 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7704 N$15408 N$15407 "Straight Waveguide" sch_x=-87 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7705 N$15410 N$15409 "Straight Waveguide" sch_x=-87 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7706 N$15412 N$15411 "Straight Waveguide" sch_x=-87 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7707 N$15414 N$15413 "Straight Waveguide" sch_x=-87 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7708 N$15416 N$15415 "Straight Waveguide" sch_x=-87 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7709 N$15418 N$15417 "Straight Waveguide" sch_x=-85 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7710 N$15420 N$15419 "Straight Waveguide" sch_x=-85 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7711 N$15422 N$15421 "Straight Waveguide" sch_x=-85 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7712 N$15424 N$15423 "Straight Waveguide" sch_x=-85 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7713 N$15426 N$15425 "Straight Waveguide" sch_x=-85 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7714 N$15428 N$15427 "Straight Waveguide" sch_x=-85 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7715 N$15430 N$15429 "Straight Waveguide" sch_x=-85 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7716 N$15432 N$15431 "Straight Waveguide" sch_x=-85 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7717 N$15434 N$15433 "Straight Waveguide" sch_x=-85 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7718 N$15436 N$15435 "Straight Waveguide" sch_x=-85 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7719 N$15438 N$15437 "Straight Waveguide" sch_x=-85 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7720 N$15440 N$15439 "Straight Waveguide" sch_x=-85 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7721 N$15442 N$15441 "Straight Waveguide" sch_x=-85 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7722 N$15444 N$15443 "Straight Waveguide" sch_x=-85 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7723 N$15446 N$15445 "Straight Waveguide" sch_x=-85 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7724 N$15448 N$15447 "Straight Waveguide" sch_x=-85 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7725 N$15450 N$15449 "Straight Waveguide" sch_x=-85 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7726 N$15452 N$15451 "Straight Waveguide" sch_x=-85 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7727 N$15454 N$15453 "Straight Waveguide" sch_x=-85 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7728 N$15456 N$15455 "Straight Waveguide" sch_x=-85 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7729 N$15458 N$15457 "Straight Waveguide" sch_x=-85 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7730 N$15460 N$15459 "Straight Waveguide" sch_x=-85 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7731 N$15462 N$15461 "Straight Waveguide" sch_x=-83 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7732 N$15464 N$15463 "Straight Waveguide" sch_x=-83 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7733 N$15466 N$15465 "Straight Waveguide" sch_x=-83 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7734 N$15468 N$15467 "Straight Waveguide" sch_x=-83 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7735 N$15470 N$15469 "Straight Waveguide" sch_x=-83 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7736 N$15472 N$15471 "Straight Waveguide" sch_x=-83 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7737 N$15474 N$15473 "Straight Waveguide" sch_x=-83 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7738 N$15476 N$15475 "Straight Waveguide" sch_x=-83 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7739 N$15478 N$15477 "Straight Waveguide" sch_x=-83 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7740 N$15480 N$15479 "Straight Waveguide" sch_x=-83 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7741 N$15482 N$15481 "Straight Waveguide" sch_x=-83 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7742 N$15484 N$15483 "Straight Waveguide" sch_x=-83 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7743 N$15486 N$15485 "Straight Waveguide" sch_x=-83 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7744 N$15488 N$15487 "Straight Waveguide" sch_x=-83 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7745 N$15490 N$15489 "Straight Waveguide" sch_x=-83 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7746 N$15492 N$15491 "Straight Waveguide" sch_x=-83 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7747 N$15494 N$15493 "Straight Waveguide" sch_x=-83 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7748 N$15496 N$15495 "Straight Waveguide" sch_x=-83 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7749 N$15498 N$15497 "Straight Waveguide" sch_x=-83 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7750 N$15500 N$15499 "Straight Waveguide" sch_x=-83 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7751 N$15502 N$15501 "Straight Waveguide" sch_x=-81 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7752 N$15504 N$15503 "Straight Waveguide" sch_x=-81 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7753 N$15506 N$15505 "Straight Waveguide" sch_x=-81 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7754 N$15508 N$15507 "Straight Waveguide" sch_x=-81 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7755 N$15510 N$15509 "Straight Waveguide" sch_x=-81 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7756 N$15512 N$15511 "Straight Waveguide" sch_x=-81 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7757 N$15514 N$15513 "Straight Waveguide" sch_x=-81 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7758 N$15516 N$15515 "Straight Waveguide" sch_x=-81 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7759 N$15518 N$15517 "Straight Waveguide" sch_x=-81 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7760 N$15520 N$15519 "Straight Waveguide" sch_x=-81 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7761 N$15522 N$15521 "Straight Waveguide" sch_x=-81 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7762 N$15524 N$15523 "Straight Waveguide" sch_x=-81 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7763 N$15526 N$15525 "Straight Waveguide" sch_x=-81 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7764 N$15528 N$15527 "Straight Waveguide" sch_x=-81 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7765 N$15530 N$15529 "Straight Waveguide" sch_x=-81 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7766 N$15532 N$15531 "Straight Waveguide" sch_x=-81 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7767 N$15534 N$15533 "Straight Waveguide" sch_x=-81 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7768 N$15536 N$15535 "Straight Waveguide" sch_x=-81 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7769 N$15538 N$15537 "Straight Waveguide" sch_x=-79 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7770 N$15540 N$15539 "Straight Waveguide" sch_x=-79 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7771 N$15542 N$15541 "Straight Waveguide" sch_x=-79 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7772 N$15544 N$15543 "Straight Waveguide" sch_x=-79 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7773 N$15546 N$15545 "Straight Waveguide" sch_x=-79 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7774 N$15548 N$15547 "Straight Waveguide" sch_x=-79 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7775 N$15550 N$15549 "Straight Waveguide" sch_x=-79 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7776 N$15552 N$15551 "Straight Waveguide" sch_x=-79 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7777 N$15554 N$15553 "Straight Waveguide" sch_x=-79 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7778 N$15556 N$15555 "Straight Waveguide" sch_x=-79 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7779 N$15558 N$15557 "Straight Waveguide" sch_x=-79 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7780 N$15560 N$15559 "Straight Waveguide" sch_x=-79 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7781 N$15562 N$15561 "Straight Waveguide" sch_x=-79 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7782 N$15564 N$15563 "Straight Waveguide" sch_x=-79 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7783 N$15566 N$15565 "Straight Waveguide" sch_x=-79 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7784 N$15568 N$15567 "Straight Waveguide" sch_x=-79 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7785 N$15570 N$15569 "Straight Waveguide" sch_x=-77 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7786 N$15572 N$15571 "Straight Waveguide" sch_x=-77 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7787 N$15574 N$15573 "Straight Waveguide" sch_x=-77 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7788 N$15576 N$15575 "Straight Waveguide" sch_x=-77 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7789 N$15578 N$15577 "Straight Waveguide" sch_x=-77 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7790 N$15580 N$15579 "Straight Waveguide" sch_x=-77 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7791 N$15582 N$15581 "Straight Waveguide" sch_x=-77 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7792 N$15584 N$15583 "Straight Waveguide" sch_x=-77 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7793 N$15586 N$15585 "Straight Waveguide" sch_x=-77 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7794 N$15588 N$15587 "Straight Waveguide" sch_x=-77 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7795 N$15590 N$15589 "Straight Waveguide" sch_x=-77 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7796 N$15592 N$15591 "Straight Waveguide" sch_x=-77 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7797 N$15594 N$15593 "Straight Waveguide" sch_x=-77 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7798 N$15596 N$15595 "Straight Waveguide" sch_x=-77 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7799 N$15598 N$15597 "Straight Waveguide" sch_x=-75 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7800 N$15600 N$15599 "Straight Waveguide" sch_x=-75 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7801 N$15602 N$15601 "Straight Waveguide" sch_x=-75 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7802 N$15604 N$15603 "Straight Waveguide" sch_x=-75 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7803 N$15606 N$15605 "Straight Waveguide" sch_x=-75 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7804 N$15608 N$15607 "Straight Waveguide" sch_x=-75 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7805 N$15610 N$15609 "Straight Waveguide" sch_x=-75 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7806 N$15612 N$15611 "Straight Waveguide" sch_x=-75 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7807 N$15614 N$15613 "Straight Waveguide" sch_x=-75 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7808 N$15616 N$15615 "Straight Waveguide" sch_x=-75 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7809 N$15618 N$15617 "Straight Waveguide" sch_x=-75 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7810 N$15620 N$15619 "Straight Waveguide" sch_x=-75 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7811 N$15622 N$15621 "Straight Waveguide" sch_x=-73 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7812 N$15624 N$15623 "Straight Waveguide" sch_x=-73 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7813 N$15626 N$15625 "Straight Waveguide" sch_x=-73 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7814 N$15628 N$15627 "Straight Waveguide" sch_x=-73 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7815 N$15630 N$15629 "Straight Waveguide" sch_x=-73 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7816 N$15632 N$15631 "Straight Waveguide" sch_x=-73 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7817 N$15634 N$15633 "Straight Waveguide" sch_x=-73 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7818 N$15636 N$15635 "Straight Waveguide" sch_x=-73 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7819 N$15638 N$15637 "Straight Waveguide" sch_x=-73 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7820 N$15640 N$15639 "Straight Waveguide" sch_x=-73 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7821 N$15642 N$15641 "Straight Waveguide" sch_x=-71 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7822 N$15644 N$15643 "Straight Waveguide" sch_x=-71 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7823 N$15646 N$15645 "Straight Waveguide" sch_x=-71 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7824 N$15648 N$15647 "Straight Waveguide" sch_x=-71 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7825 N$15650 N$15649 "Straight Waveguide" sch_x=-71 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7826 N$15652 N$15651 "Straight Waveguide" sch_x=-71 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7827 N$15654 N$15653 "Straight Waveguide" sch_x=-71 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7828 N$15656 N$15655 "Straight Waveguide" sch_x=-71 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7829 N$15658 N$15657 "Straight Waveguide" sch_x=-69 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7830 N$15660 N$15659 "Straight Waveguide" sch_x=-69 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7831 N$15662 N$15661 "Straight Waveguide" sch_x=-69 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7832 N$15664 N$15663 "Straight Waveguide" sch_x=-69 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7833 N$15666 N$15665 "Straight Waveguide" sch_x=-69 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7834 N$15668 N$15667 "Straight Waveguide" sch_x=-69 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7835 N$15670 N$15669 "Straight Waveguide" sch_x=-67 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7836 N$15672 N$15671 "Straight Waveguide" sch_x=-67 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7837 N$15674 N$15673 "Straight Waveguide" sch_x=-67 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7838 N$15676 N$15675 "Straight Waveguide" sch_x=-67 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7839 N$15678 N$15677 "Straight Waveguide" sch_x=-65 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7840 N$15680 N$15679 "Straight Waveguide" sch_x=-65 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7841 N$15681 N$15682 "Straight Waveguide" sch_x=-93 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7842 N$15683 N$15684 "Straight Waveguide" sch_x=-92 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7843 N$15685 N$15686 "Straight Waveguide" sch_x=-91 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7844 N$15687 N$15688 "Straight Waveguide" sch_x=-90 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7845 N$15689 N$15690 "Straight Waveguide" sch_x=-89 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7846 N$15691 N$15692 "Straight Waveguide" sch_x=-88 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7847 N$15693 N$15694 "Straight Waveguide" sch_x=-87 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7848 N$15695 N$15696 "Straight Waveguide" sch_x=-86 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7849 N$15697 N$15698 "Straight Waveguide" sch_x=-85 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7850 N$15699 N$15700 "Straight Waveguide" sch_x=-84 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7851 N$15701 N$15702 "Straight Waveguide" sch_x=-83 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7852 N$15703 N$15704 "Straight Waveguide" sch_x=-82 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7853 N$15705 N$15706 "Straight Waveguide" sch_x=-81 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7854 N$15707 N$15708 "Straight Waveguide" sch_x=-80 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7855 N$15709 N$15710 "Straight Waveguide" sch_x=-79 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7856 N$15711 N$15712 "Straight Waveguide" sch_x=-78 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7857 N$15713 N$15714 "Straight Waveguide" sch_x=-77 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7858 N$15715 N$15716 "Straight Waveguide" sch_x=-76 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7859 N$15717 N$15718 "Straight Waveguide" sch_x=-75 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7860 N$15719 N$15720 "Straight Waveguide" sch_x=-74 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7861 N$15721 N$15722 "Straight Waveguide" sch_x=-73 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7862 N$15723 N$15724 "Straight Waveguide" sch_x=-72 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7863 N$15725 N$15726 "Straight Waveguide" sch_x=-71 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7864 N$15727 N$15728 "Straight Waveguide" sch_x=-70 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7865 N$15729 N$15730 "Straight Waveguide" sch_x=-69 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7866 N$15731 N$15732 "Straight Waveguide" sch_x=-68 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7867 N$15733 N$15734 "Straight Waveguide" sch_x=-67 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7868 N$15735 N$15736 "Straight Waveguide" sch_x=-66 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7869 N$15737 N$15738 "Straight Waveguide" sch_x=-65 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7870 N$15739 N$15740 "Straight Waveguide" sch_x=-64 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7871 N$15741 N$15742 "Straight Waveguide" sch_x=-63 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7872 N$15743 N$15744 "Straight Waveguide" sch_x=-63 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7873 N$15745 N$15746 "Straight Waveguide" sch_x=-64 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7874 N$15747 N$15748 "Straight Waveguide" sch_x=-65 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7875 N$15749 N$15750 "Straight Waveguide" sch_x=-66 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7876 N$15751 N$15752 "Straight Waveguide" sch_x=-67 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7877 N$15753 N$15754 "Straight Waveguide" sch_x=-68 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7878 N$15755 N$15756 "Straight Waveguide" sch_x=-69 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7879 N$15757 N$15758 "Straight Waveguide" sch_x=-70 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7880 N$15759 N$15760 "Straight Waveguide" sch_x=-71 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7881 N$15761 N$15762 "Straight Waveguide" sch_x=-72 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7882 N$15763 N$15764 "Straight Waveguide" sch_x=-73 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7883 N$15765 N$15766 "Straight Waveguide" sch_x=-74 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7884 N$15767 N$15768 "Straight Waveguide" sch_x=-75 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7885 N$15769 N$15770 "Straight Waveguide" sch_x=-76 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7886 N$15771 N$15772 "Straight Waveguide" sch_x=-77 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7887 N$15773 N$15774 "Straight Waveguide" sch_x=-78 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7888 N$15775 N$15776 "Straight Waveguide" sch_x=-79 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7889 N$15777 N$15778 "Straight Waveguide" sch_x=-80 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7890 N$15779 N$15780 "Straight Waveguide" sch_x=-81 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7891 N$15781 N$15782 "Straight Waveguide" sch_x=-82 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7892 N$15783 N$15784 "Straight Waveguide" sch_x=-83 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7893 N$15785 N$15786 "Straight Waveguide" sch_x=-84 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7894 N$15787 N$15788 "Straight Waveguide" sch_x=-85 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7895 N$15789 N$15790 "Straight Waveguide" sch_x=-86 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7896 N$15791 N$15792 "Straight Waveguide" sch_x=-87 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7897 N$15793 N$15794 "Straight Waveguide" sch_x=-88 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7898 N$15795 N$15796 "Straight Waveguide" sch_x=-89 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7899 N$15797 N$15798 "Straight Waveguide" sch_x=-90 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7900 N$15799 N$15800 "Straight Waveguide" sch_x=-91 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7901 N$15801 N$15802 "Straight Waveguide" sch_x=-92 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7902 N$15803 N$15804 "Straight Waveguide" sch_x=-93 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7903 N$15805 N$15806 "Straight Waveguide" sch_x=-94 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7904 N$15807 N$15808 "Straight Waveguide" sch_x=-94 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7905 N$15809 N$15810 "Straight Waveguide" sch_x=125 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7906 N$15811 N$15812 "Straight Waveguide" sch_x=125 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7907 N$15813 N$15814 "Straight Waveguide" sch_x=125 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7908 N$15815 N$15816 "Straight Waveguide" sch_x=125 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7909 N$15817 N$15818 "Straight Waveguide" sch_x=125 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7910 N$15819 N$15820 "Straight Waveguide" sch_x=125 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7911 N$15821 N$15822 "Straight Waveguide" sch_x=125 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7912 N$15823 N$15824 "Straight Waveguide" sch_x=125 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7913 N$15825 N$15826 "Straight Waveguide" sch_x=125 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7914 N$15827 N$15828 "Straight Waveguide" sch_x=125 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7915 N$15829 N$15830 "Straight Waveguide" sch_x=125 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7916 N$15831 N$15832 "Straight Waveguide" sch_x=125 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7917 N$15833 N$15834 "Straight Waveguide" sch_x=125 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7918 N$15835 N$15836 "Straight Waveguide" sch_x=125 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7919 N$15837 N$15838 "Straight Waveguide" sch_x=125 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7920 N$15839 N$15840 "Straight Waveguide" sch_x=125 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7921 N$15841 N$15842 "Straight Waveguide" sch_x=125 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7922 N$15843 N$15844 "Straight Waveguide" sch_x=125 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7923 N$15845 N$15846 "Straight Waveguide" sch_x=125 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7924 N$15847 N$15848 "Straight Waveguide" sch_x=125 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7925 N$15849 N$15850 "Straight Waveguide" sch_x=125 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7926 N$15851 N$15852 "Straight Waveguide" sch_x=125 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7927 N$15853 N$15854 "Straight Waveguide" sch_x=125 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7928 N$15855 N$15856 "Straight Waveguide" sch_x=125 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7929 N$15857 N$15858 "Straight Waveguide" sch_x=125 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7930 N$15859 N$15860 "Straight Waveguide" sch_x=125 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7931 N$15861 N$15862 "Straight Waveguide" sch_x=125 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7932 N$15863 N$15864 "Straight Waveguide" sch_x=125 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7933 N$15865 N$15866 "Straight Waveguide" sch_x=125 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7934 N$15867 N$15868 "Straight Waveguide" sch_x=125 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7935 N$15869 N$15870 "Straight Waveguide" sch_x=125 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7936 N$15871 N$15872 "Straight Waveguide" sch_x=125 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7937 N$15873 N$15874 "Straight Waveguide" sch_x=125 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7938 N$15875 N$15876 "Straight Waveguide" sch_x=125 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7939 N$15877 N$15878 "Straight Waveguide" sch_x=125 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7940 N$15879 N$15880 "Straight Waveguide" sch_x=125 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7941 N$15881 N$15882 "Straight Waveguide" sch_x=125 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7942 N$15883 N$15884 "Straight Waveguide" sch_x=125 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7943 N$15885 N$15886 "Straight Waveguide" sch_x=125 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7944 N$15887 N$15888 "Straight Waveguide" sch_x=125 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7945 N$15889 N$15890 "Straight Waveguide" sch_x=125 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7946 N$15891 N$15892 "Straight Waveguide" sch_x=125 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7947 N$15893 N$15894 "Straight Waveguide" sch_x=125 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7948 N$15895 N$15896 "Straight Waveguide" sch_x=125 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7949 N$15897 N$15898 "Straight Waveguide" sch_x=125 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7950 N$15899 N$15900 "Straight Waveguide" sch_x=125 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7951 N$15901 N$15902 "Straight Waveguide" sch_x=125 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7952 N$15903 N$15904 "Straight Waveguide" sch_x=125 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7953 N$15905 N$15906 "Straight Waveguide" sch_x=125 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7954 N$15907 N$15908 "Straight Waveguide" sch_x=125 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7955 N$15909 N$15910 "Straight Waveguide" sch_x=125 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7956 N$15911 N$15912 "Straight Waveguide" sch_x=125 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7957 N$15913 N$15914 "Straight Waveguide" sch_x=125 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7958 N$15915 N$15916 "Straight Waveguide" sch_x=125 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7959 N$15917 N$15918 "Straight Waveguide" sch_x=125 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7960 N$15919 N$15920 "Straight Waveguide" sch_x=125 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7961 N$15921 N$15922 "Straight Waveguide" sch_x=125 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7962 N$15923 N$15924 "Straight Waveguide" sch_x=125 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7963 N$15925 N$15926 "Straight Waveguide" sch_x=125 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7964 N$15927 N$15928 "Straight Waveguide" sch_x=125 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7965 N$15929 N$15930 "Straight Waveguide" sch_x=125 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7966 N$15931 N$15932 "Straight Waveguide" sch_x=125 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7967 N$15933 N$15934 "Straight Waveguide" sch_x=123 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7968 N$15935 N$15936 "Straight Waveguide" sch_x=123 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7969 N$15937 N$15938 "Straight Waveguide" sch_x=123 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7970 N$15939 N$15940 "Straight Waveguide" sch_x=123 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7971 N$15941 N$15942 "Straight Waveguide" sch_x=123 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7972 N$15943 N$15944 "Straight Waveguide" sch_x=123 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7973 N$15945 N$15946 "Straight Waveguide" sch_x=123 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7974 N$15947 N$15948 "Straight Waveguide" sch_x=123 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7975 N$15949 N$15950 "Straight Waveguide" sch_x=123 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7976 N$15951 N$15952 "Straight Waveguide" sch_x=123 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7977 N$15953 N$15954 "Straight Waveguide" sch_x=123 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7978 N$15955 N$15956 "Straight Waveguide" sch_x=123 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7979 N$15957 N$15958 "Straight Waveguide" sch_x=123 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7980 N$15959 N$15960 "Straight Waveguide" sch_x=123 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7981 N$15961 N$15962 "Straight Waveguide" sch_x=123 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7982 N$15963 N$15964 "Straight Waveguide" sch_x=123 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7983 N$15965 N$15966 "Straight Waveguide" sch_x=123 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7984 N$15967 N$15968 "Straight Waveguide" sch_x=123 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7985 N$15969 N$15970 "Straight Waveguide" sch_x=123 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7986 N$15971 N$15972 "Straight Waveguide" sch_x=123 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7987 N$15973 N$15974 "Straight Waveguide" sch_x=123 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7988 N$15975 N$15976 "Straight Waveguide" sch_x=123 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7989 N$15977 N$15978 "Straight Waveguide" sch_x=123 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7990 N$15979 N$15980 "Straight Waveguide" sch_x=123 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7991 N$15981 N$15982 "Straight Waveguide" sch_x=123 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7992 N$15983 N$15984 "Straight Waveguide" sch_x=123 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7993 N$15985 N$15986 "Straight Waveguide" sch_x=123 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7994 N$15987 N$15988 "Straight Waveguide" sch_x=123 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7995 N$15989 N$15990 "Straight Waveguide" sch_x=123 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7996 N$15991 N$15992 "Straight Waveguide" sch_x=123 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7997 N$15993 N$15994 "Straight Waveguide" sch_x=123 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7998 N$15995 N$15996 "Straight Waveguide" sch_x=123 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7999 N$15997 N$15998 "Straight Waveguide" sch_x=123 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8000 N$15999 N$16000 "Straight Waveguide" sch_x=123 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8001 N$16001 N$16002 "Straight Waveguide" sch_x=123 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8002 N$16003 N$16004 "Straight Waveguide" sch_x=123 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8003 N$16005 N$16006 "Straight Waveguide" sch_x=123 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8004 N$16007 N$16008 "Straight Waveguide" sch_x=123 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8005 N$16009 N$16010 "Straight Waveguide" sch_x=123 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8006 N$16011 N$16012 "Straight Waveguide" sch_x=123 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8007 N$16013 N$16014 "Straight Waveguide" sch_x=123 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8008 N$16015 N$16016 "Straight Waveguide" sch_x=123 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8009 N$16017 N$16018 "Straight Waveguide" sch_x=123 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8010 N$16019 N$16020 "Straight Waveguide" sch_x=123 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8011 N$16021 N$16022 "Straight Waveguide" sch_x=123 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8012 N$16023 N$16024 "Straight Waveguide" sch_x=123 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8013 N$16025 N$16026 "Straight Waveguide" sch_x=123 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8014 N$16027 N$16028 "Straight Waveguide" sch_x=123 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8015 N$16029 N$16030 "Straight Waveguide" sch_x=123 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8016 N$16031 N$16032 "Straight Waveguide" sch_x=123 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8017 N$16033 N$16034 "Straight Waveguide" sch_x=123 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8018 N$16035 N$16036 "Straight Waveguide" sch_x=123 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8019 N$16037 N$16038 "Straight Waveguide" sch_x=123 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8020 N$16039 N$16040 "Straight Waveguide" sch_x=123 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8021 N$16041 N$16042 "Straight Waveguide" sch_x=123 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8022 N$16043 N$16044 "Straight Waveguide" sch_x=123 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8023 N$16045 N$16046 "Straight Waveguide" sch_x=123 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8024 N$16047 N$16048 "Straight Waveguide" sch_x=123 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8025 N$16049 N$16050 "Straight Waveguide" sch_x=123 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8026 N$16051 N$16052 "Straight Waveguide" sch_x=123 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8027 N$16053 N$16054 "Straight Waveguide" sch_x=121 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8028 N$16055 N$16056 "Straight Waveguide" sch_x=121 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8029 N$16057 N$16058 "Straight Waveguide" sch_x=121 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8030 N$16059 N$16060 "Straight Waveguide" sch_x=121 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8031 N$16061 N$16062 "Straight Waveguide" sch_x=121 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8032 N$16063 N$16064 "Straight Waveguide" sch_x=121 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8033 N$16065 N$16066 "Straight Waveguide" sch_x=121 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8034 N$16067 N$16068 "Straight Waveguide" sch_x=121 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8035 N$16069 N$16070 "Straight Waveguide" sch_x=121 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8036 N$16071 N$16072 "Straight Waveguide" sch_x=121 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8037 N$16073 N$16074 "Straight Waveguide" sch_x=121 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8038 N$16075 N$16076 "Straight Waveguide" sch_x=121 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8039 N$16077 N$16078 "Straight Waveguide" sch_x=121 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8040 N$16079 N$16080 "Straight Waveguide" sch_x=121 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8041 N$16081 N$16082 "Straight Waveguide" sch_x=121 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8042 N$16083 N$16084 "Straight Waveguide" sch_x=121 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8043 N$16085 N$16086 "Straight Waveguide" sch_x=121 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8044 N$16087 N$16088 "Straight Waveguide" sch_x=121 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8045 N$16089 N$16090 "Straight Waveguide" sch_x=121 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8046 N$16091 N$16092 "Straight Waveguide" sch_x=121 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8047 N$16093 N$16094 "Straight Waveguide" sch_x=121 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8048 N$16095 N$16096 "Straight Waveguide" sch_x=121 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8049 N$16097 N$16098 "Straight Waveguide" sch_x=121 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8050 N$16099 N$16100 "Straight Waveguide" sch_x=121 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8051 N$16101 N$16102 "Straight Waveguide" sch_x=121 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8052 N$16103 N$16104 "Straight Waveguide" sch_x=121 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8053 N$16105 N$16106 "Straight Waveguide" sch_x=121 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8054 N$16107 N$16108 "Straight Waveguide" sch_x=121 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8055 N$16109 N$16110 "Straight Waveguide" sch_x=121 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8056 N$16111 N$16112 "Straight Waveguide" sch_x=121 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8057 N$16113 N$16114 "Straight Waveguide" sch_x=121 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8058 N$16115 N$16116 "Straight Waveguide" sch_x=121 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8059 N$16117 N$16118 "Straight Waveguide" sch_x=121 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8060 N$16119 N$16120 "Straight Waveguide" sch_x=121 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8061 N$16121 N$16122 "Straight Waveguide" sch_x=121 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8062 N$16123 N$16124 "Straight Waveguide" sch_x=121 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8063 N$16125 N$16126 "Straight Waveguide" sch_x=121 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8064 N$16127 N$16128 "Straight Waveguide" sch_x=121 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8065 N$16129 N$16130 "Straight Waveguide" sch_x=121 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8066 N$16131 N$16132 "Straight Waveguide" sch_x=121 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8067 N$16133 N$16134 "Straight Waveguide" sch_x=121 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8068 N$16135 N$16136 "Straight Waveguide" sch_x=121 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8069 N$16137 N$16138 "Straight Waveguide" sch_x=121 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8070 N$16139 N$16140 "Straight Waveguide" sch_x=121 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8071 N$16141 N$16142 "Straight Waveguide" sch_x=121 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8072 N$16143 N$16144 "Straight Waveguide" sch_x=121 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8073 N$16145 N$16146 "Straight Waveguide" sch_x=121 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8074 N$16147 N$16148 "Straight Waveguide" sch_x=121 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8075 N$16149 N$16150 "Straight Waveguide" sch_x=121 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8076 N$16151 N$16152 "Straight Waveguide" sch_x=121 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8077 N$16153 N$16154 "Straight Waveguide" sch_x=121 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8078 N$16155 N$16156 "Straight Waveguide" sch_x=121 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8079 N$16157 N$16158 "Straight Waveguide" sch_x=121 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8080 N$16159 N$16160 "Straight Waveguide" sch_x=121 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8081 N$16161 N$16162 "Straight Waveguide" sch_x=121 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8082 N$16163 N$16164 "Straight Waveguide" sch_x=121 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8083 N$16165 N$16166 "Straight Waveguide" sch_x=121 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8084 N$16167 N$16168 "Straight Waveguide" sch_x=121 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8085 N$16169 N$16170 "Straight Waveguide" sch_x=119 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8086 N$16171 N$16172 "Straight Waveguide" sch_x=119 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8087 N$16173 N$16174 "Straight Waveguide" sch_x=119 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8088 N$16175 N$16176 "Straight Waveguide" sch_x=119 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8089 N$16177 N$16178 "Straight Waveguide" sch_x=119 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8090 N$16179 N$16180 "Straight Waveguide" sch_x=119 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8091 N$16181 N$16182 "Straight Waveguide" sch_x=119 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8092 N$16183 N$16184 "Straight Waveguide" sch_x=119 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8093 N$16185 N$16186 "Straight Waveguide" sch_x=119 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8094 N$16187 N$16188 "Straight Waveguide" sch_x=119 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8095 N$16189 N$16190 "Straight Waveguide" sch_x=119 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8096 N$16191 N$16192 "Straight Waveguide" sch_x=119 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8097 N$16193 N$16194 "Straight Waveguide" sch_x=119 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8098 N$16195 N$16196 "Straight Waveguide" sch_x=119 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8099 N$16197 N$16198 "Straight Waveguide" sch_x=119 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8100 N$16199 N$16200 "Straight Waveguide" sch_x=119 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8101 N$16201 N$16202 "Straight Waveguide" sch_x=119 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8102 N$16203 N$16204 "Straight Waveguide" sch_x=119 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8103 N$16205 N$16206 "Straight Waveguide" sch_x=119 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8104 N$16207 N$16208 "Straight Waveguide" sch_x=119 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8105 N$16209 N$16210 "Straight Waveguide" sch_x=119 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8106 N$16211 N$16212 "Straight Waveguide" sch_x=119 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8107 N$16213 N$16214 "Straight Waveguide" sch_x=119 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8108 N$16215 N$16216 "Straight Waveguide" sch_x=119 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8109 N$16217 N$16218 "Straight Waveguide" sch_x=119 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8110 N$16219 N$16220 "Straight Waveguide" sch_x=119 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8111 N$16221 N$16222 "Straight Waveguide" sch_x=119 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8112 N$16223 N$16224 "Straight Waveguide" sch_x=119 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8113 N$16225 N$16226 "Straight Waveguide" sch_x=119 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8114 N$16227 N$16228 "Straight Waveguide" sch_x=119 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8115 N$16229 N$16230 "Straight Waveguide" sch_x=119 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8116 N$16231 N$16232 "Straight Waveguide" sch_x=119 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8117 N$16233 N$16234 "Straight Waveguide" sch_x=119 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8118 N$16235 N$16236 "Straight Waveguide" sch_x=119 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8119 N$16237 N$16238 "Straight Waveguide" sch_x=119 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8120 N$16239 N$16240 "Straight Waveguide" sch_x=119 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8121 N$16241 N$16242 "Straight Waveguide" sch_x=119 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8122 N$16243 N$16244 "Straight Waveguide" sch_x=119 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8123 N$16245 N$16246 "Straight Waveguide" sch_x=119 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8124 N$16247 N$16248 "Straight Waveguide" sch_x=119 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8125 N$16249 N$16250 "Straight Waveguide" sch_x=119 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8126 N$16251 N$16252 "Straight Waveguide" sch_x=119 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8127 N$16253 N$16254 "Straight Waveguide" sch_x=119 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8128 N$16255 N$16256 "Straight Waveguide" sch_x=119 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8129 N$16257 N$16258 "Straight Waveguide" sch_x=119 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8130 N$16259 N$16260 "Straight Waveguide" sch_x=119 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8131 N$16261 N$16262 "Straight Waveguide" sch_x=119 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8132 N$16263 N$16264 "Straight Waveguide" sch_x=119 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8133 N$16265 N$16266 "Straight Waveguide" sch_x=119 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8134 N$16267 N$16268 "Straight Waveguide" sch_x=119 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8135 N$16269 N$16270 "Straight Waveguide" sch_x=119 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8136 N$16271 N$16272 "Straight Waveguide" sch_x=119 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8137 N$16273 N$16274 "Straight Waveguide" sch_x=119 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8138 N$16275 N$16276 "Straight Waveguide" sch_x=119 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8139 N$16277 N$16278 "Straight Waveguide" sch_x=119 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8140 N$16279 N$16280 "Straight Waveguide" sch_x=119 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8141 N$16281 N$16282 "Straight Waveguide" sch_x=117 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8142 N$16283 N$16284 "Straight Waveguide" sch_x=117 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8143 N$16285 N$16286 "Straight Waveguide" sch_x=117 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8144 N$16287 N$16288 "Straight Waveguide" sch_x=117 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8145 N$16289 N$16290 "Straight Waveguide" sch_x=117 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8146 N$16291 N$16292 "Straight Waveguide" sch_x=117 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8147 N$16293 N$16294 "Straight Waveguide" sch_x=117 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8148 N$16295 N$16296 "Straight Waveguide" sch_x=117 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8149 N$16297 N$16298 "Straight Waveguide" sch_x=117 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8150 N$16299 N$16300 "Straight Waveguide" sch_x=117 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8151 N$16301 N$16302 "Straight Waveguide" sch_x=117 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8152 N$16303 N$16304 "Straight Waveguide" sch_x=117 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8153 N$16305 N$16306 "Straight Waveguide" sch_x=117 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8154 N$16307 N$16308 "Straight Waveguide" sch_x=117 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8155 N$16309 N$16310 "Straight Waveguide" sch_x=117 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8156 N$16311 N$16312 "Straight Waveguide" sch_x=117 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8157 N$16313 N$16314 "Straight Waveguide" sch_x=117 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8158 N$16315 N$16316 "Straight Waveguide" sch_x=117 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8159 N$16317 N$16318 "Straight Waveguide" sch_x=117 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8160 N$16319 N$16320 "Straight Waveguide" sch_x=117 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8161 N$16321 N$16322 "Straight Waveguide" sch_x=117 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8162 N$16323 N$16324 "Straight Waveguide" sch_x=117 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8163 N$16325 N$16326 "Straight Waveguide" sch_x=117 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8164 N$16327 N$16328 "Straight Waveguide" sch_x=117 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8165 N$16329 N$16330 "Straight Waveguide" sch_x=117 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8166 N$16331 N$16332 "Straight Waveguide" sch_x=117 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8167 N$16333 N$16334 "Straight Waveguide" sch_x=117 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8168 N$16335 N$16336 "Straight Waveguide" sch_x=117 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8169 N$16337 N$16338 "Straight Waveguide" sch_x=117 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8170 N$16339 N$16340 "Straight Waveguide" sch_x=117 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8171 N$16341 N$16342 "Straight Waveguide" sch_x=117 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8172 N$16343 N$16344 "Straight Waveguide" sch_x=117 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8173 N$16345 N$16346 "Straight Waveguide" sch_x=117 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8174 N$16347 N$16348 "Straight Waveguide" sch_x=117 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8175 N$16349 N$16350 "Straight Waveguide" sch_x=117 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8176 N$16351 N$16352 "Straight Waveguide" sch_x=117 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8177 N$16353 N$16354 "Straight Waveguide" sch_x=117 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8178 N$16355 N$16356 "Straight Waveguide" sch_x=117 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8179 N$16357 N$16358 "Straight Waveguide" sch_x=117 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8180 N$16359 N$16360 "Straight Waveguide" sch_x=117 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8181 N$16361 N$16362 "Straight Waveguide" sch_x=117 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8182 N$16363 N$16364 "Straight Waveguide" sch_x=117 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8183 N$16365 N$16366 "Straight Waveguide" sch_x=117 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8184 N$16367 N$16368 "Straight Waveguide" sch_x=117 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8185 N$16369 N$16370 "Straight Waveguide" sch_x=117 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8186 N$16371 N$16372 "Straight Waveguide" sch_x=117 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8187 N$16373 N$16374 "Straight Waveguide" sch_x=117 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8188 N$16375 N$16376 "Straight Waveguide" sch_x=117 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8189 N$16377 N$16378 "Straight Waveguide" sch_x=117 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8190 N$16379 N$16380 "Straight Waveguide" sch_x=117 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8191 N$16381 N$16382 "Straight Waveguide" sch_x=117 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8192 N$16383 N$16384 "Straight Waveguide" sch_x=117 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8193 N$16385 N$16386 "Straight Waveguide" sch_x=117 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8194 N$16387 N$16388 "Straight Waveguide" sch_x=117 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8195 N$16389 N$16390 "Straight Waveguide" sch_x=115 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8196 N$16391 N$16392 "Straight Waveguide" sch_x=115 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8197 N$16393 N$16394 "Straight Waveguide" sch_x=115 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8198 N$16395 N$16396 "Straight Waveguide" sch_x=115 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8199 N$16397 N$16398 "Straight Waveguide" sch_x=115 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8200 N$16399 N$16400 "Straight Waveguide" sch_x=115 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8201 N$16401 N$16402 "Straight Waveguide" sch_x=115 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8202 N$16403 N$16404 "Straight Waveguide" sch_x=115 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8203 N$16405 N$16406 "Straight Waveguide" sch_x=115 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8204 N$16407 N$16408 "Straight Waveguide" sch_x=115 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8205 N$16409 N$16410 "Straight Waveguide" sch_x=115 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8206 N$16411 N$16412 "Straight Waveguide" sch_x=115 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8207 N$16413 N$16414 "Straight Waveguide" sch_x=115 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8208 N$16415 N$16416 "Straight Waveguide" sch_x=115 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8209 N$16417 N$16418 "Straight Waveguide" sch_x=115 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8210 N$16419 N$16420 "Straight Waveguide" sch_x=115 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8211 N$16421 N$16422 "Straight Waveguide" sch_x=115 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8212 N$16423 N$16424 "Straight Waveguide" sch_x=115 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8213 N$16425 N$16426 "Straight Waveguide" sch_x=115 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8214 N$16427 N$16428 "Straight Waveguide" sch_x=115 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8215 N$16429 N$16430 "Straight Waveguide" sch_x=115 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8216 N$16431 N$16432 "Straight Waveguide" sch_x=115 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8217 N$16433 N$16434 "Straight Waveguide" sch_x=115 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8218 N$16435 N$16436 "Straight Waveguide" sch_x=115 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8219 N$16437 N$16438 "Straight Waveguide" sch_x=115 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8220 N$16439 N$16440 "Straight Waveguide" sch_x=115 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8221 N$16441 N$16442 "Straight Waveguide" sch_x=115 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8222 N$16443 N$16444 "Straight Waveguide" sch_x=115 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8223 N$16445 N$16446 "Straight Waveguide" sch_x=115 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8224 N$16447 N$16448 "Straight Waveguide" sch_x=115 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8225 N$16449 N$16450 "Straight Waveguide" sch_x=115 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8226 N$16451 N$16452 "Straight Waveguide" sch_x=115 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8227 N$16453 N$16454 "Straight Waveguide" sch_x=115 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8228 N$16455 N$16456 "Straight Waveguide" sch_x=115 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8229 N$16457 N$16458 "Straight Waveguide" sch_x=115 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8230 N$16459 N$16460 "Straight Waveguide" sch_x=115 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8231 N$16461 N$16462 "Straight Waveguide" sch_x=115 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8232 N$16463 N$16464 "Straight Waveguide" sch_x=115 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8233 N$16465 N$16466 "Straight Waveguide" sch_x=115 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8234 N$16467 N$16468 "Straight Waveguide" sch_x=115 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8235 N$16469 N$16470 "Straight Waveguide" sch_x=115 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8236 N$16471 N$16472 "Straight Waveguide" sch_x=115 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8237 N$16473 N$16474 "Straight Waveguide" sch_x=115 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8238 N$16475 N$16476 "Straight Waveguide" sch_x=115 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8239 N$16477 N$16478 "Straight Waveguide" sch_x=115 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8240 N$16479 N$16480 "Straight Waveguide" sch_x=115 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8241 N$16481 N$16482 "Straight Waveguide" sch_x=115 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8242 N$16483 N$16484 "Straight Waveguide" sch_x=115 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8243 N$16485 N$16486 "Straight Waveguide" sch_x=115 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8244 N$16487 N$16488 "Straight Waveguide" sch_x=115 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8245 N$16489 N$16490 "Straight Waveguide" sch_x=115 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8246 N$16491 N$16492 "Straight Waveguide" sch_x=115 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8247 N$16493 N$16494 "Straight Waveguide" sch_x=113 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8248 N$16495 N$16496 "Straight Waveguide" sch_x=113 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8249 N$16497 N$16498 "Straight Waveguide" sch_x=113 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8250 N$16499 N$16500 "Straight Waveguide" sch_x=113 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8251 N$16501 N$16502 "Straight Waveguide" sch_x=113 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8252 N$16503 N$16504 "Straight Waveguide" sch_x=113 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8253 N$16505 N$16506 "Straight Waveguide" sch_x=113 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8254 N$16507 N$16508 "Straight Waveguide" sch_x=113 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8255 N$16509 N$16510 "Straight Waveguide" sch_x=113 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8256 N$16511 N$16512 "Straight Waveguide" sch_x=113 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8257 N$16513 N$16514 "Straight Waveguide" sch_x=113 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8258 N$16515 N$16516 "Straight Waveguide" sch_x=113 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8259 N$16517 N$16518 "Straight Waveguide" sch_x=113 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8260 N$16519 N$16520 "Straight Waveguide" sch_x=113 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8261 N$16521 N$16522 "Straight Waveguide" sch_x=113 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8262 N$16523 N$16524 "Straight Waveguide" sch_x=113 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8263 N$16525 N$16526 "Straight Waveguide" sch_x=113 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8264 N$16527 N$16528 "Straight Waveguide" sch_x=113 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8265 N$16529 N$16530 "Straight Waveguide" sch_x=113 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8266 N$16531 N$16532 "Straight Waveguide" sch_x=113 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8267 N$16533 N$16534 "Straight Waveguide" sch_x=113 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8268 N$16535 N$16536 "Straight Waveguide" sch_x=113 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8269 N$16537 N$16538 "Straight Waveguide" sch_x=113 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8270 N$16539 N$16540 "Straight Waveguide" sch_x=113 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8271 N$16541 N$16542 "Straight Waveguide" sch_x=113 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8272 N$16543 N$16544 "Straight Waveguide" sch_x=113 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8273 N$16545 N$16546 "Straight Waveguide" sch_x=113 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8274 N$16547 N$16548 "Straight Waveguide" sch_x=113 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8275 N$16549 N$16550 "Straight Waveguide" sch_x=113 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8276 N$16551 N$16552 "Straight Waveguide" sch_x=113 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8277 N$16553 N$16554 "Straight Waveguide" sch_x=113 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8278 N$16555 N$16556 "Straight Waveguide" sch_x=113 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8279 N$16557 N$16558 "Straight Waveguide" sch_x=113 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8280 N$16559 N$16560 "Straight Waveguide" sch_x=113 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8281 N$16561 N$16562 "Straight Waveguide" sch_x=113 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8282 N$16563 N$16564 "Straight Waveguide" sch_x=113 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8283 N$16565 N$16566 "Straight Waveguide" sch_x=113 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8284 N$16567 N$16568 "Straight Waveguide" sch_x=113 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8285 N$16569 N$16570 "Straight Waveguide" sch_x=113 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8286 N$16571 N$16572 "Straight Waveguide" sch_x=113 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8287 N$16573 N$16574 "Straight Waveguide" sch_x=113 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8288 N$16575 N$16576 "Straight Waveguide" sch_x=113 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8289 N$16577 N$16578 "Straight Waveguide" sch_x=113 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8290 N$16579 N$16580 "Straight Waveguide" sch_x=113 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8291 N$16581 N$16582 "Straight Waveguide" sch_x=113 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8292 N$16583 N$16584 "Straight Waveguide" sch_x=113 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8293 N$16585 N$16586 "Straight Waveguide" sch_x=113 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8294 N$16587 N$16588 "Straight Waveguide" sch_x=113 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8295 N$16589 N$16590 "Straight Waveguide" sch_x=113 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8296 N$16591 N$16592 "Straight Waveguide" sch_x=113 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8297 N$16593 N$16594 "Straight Waveguide" sch_x=111 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8298 N$16595 N$16596 "Straight Waveguide" sch_x=111 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8299 N$16597 N$16598 "Straight Waveguide" sch_x=111 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8300 N$16599 N$16600 "Straight Waveguide" sch_x=111 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8301 N$16601 N$16602 "Straight Waveguide" sch_x=111 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8302 N$16603 N$16604 "Straight Waveguide" sch_x=111 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8303 N$16605 N$16606 "Straight Waveguide" sch_x=111 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8304 N$16607 N$16608 "Straight Waveguide" sch_x=111 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8305 N$16609 N$16610 "Straight Waveguide" sch_x=111 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8306 N$16611 N$16612 "Straight Waveguide" sch_x=111 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8307 N$16613 N$16614 "Straight Waveguide" sch_x=111 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8308 N$16615 N$16616 "Straight Waveguide" sch_x=111 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8309 N$16617 N$16618 "Straight Waveguide" sch_x=111 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8310 N$16619 N$16620 "Straight Waveguide" sch_x=111 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8311 N$16621 N$16622 "Straight Waveguide" sch_x=111 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8312 N$16623 N$16624 "Straight Waveguide" sch_x=111 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8313 N$16625 N$16626 "Straight Waveguide" sch_x=111 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8314 N$16627 N$16628 "Straight Waveguide" sch_x=111 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8315 N$16629 N$16630 "Straight Waveguide" sch_x=111 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8316 N$16631 N$16632 "Straight Waveguide" sch_x=111 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8317 N$16633 N$16634 "Straight Waveguide" sch_x=111 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8318 N$16635 N$16636 "Straight Waveguide" sch_x=111 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8319 N$16637 N$16638 "Straight Waveguide" sch_x=111 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8320 N$16639 N$16640 "Straight Waveguide" sch_x=111 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8321 N$16641 N$16642 "Straight Waveguide" sch_x=111 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8322 N$16643 N$16644 "Straight Waveguide" sch_x=111 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8323 N$16645 N$16646 "Straight Waveguide" sch_x=111 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8324 N$16647 N$16648 "Straight Waveguide" sch_x=111 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8325 N$16649 N$16650 "Straight Waveguide" sch_x=111 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8326 N$16651 N$16652 "Straight Waveguide" sch_x=111 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8327 N$16653 N$16654 "Straight Waveguide" sch_x=111 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8328 N$16655 N$16656 "Straight Waveguide" sch_x=111 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8329 N$16657 N$16658 "Straight Waveguide" sch_x=111 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8330 N$16659 N$16660 "Straight Waveguide" sch_x=111 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8331 N$16661 N$16662 "Straight Waveguide" sch_x=111 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8332 N$16663 N$16664 "Straight Waveguide" sch_x=111 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8333 N$16665 N$16666 "Straight Waveguide" sch_x=111 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8334 N$16667 N$16668 "Straight Waveguide" sch_x=111 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8335 N$16669 N$16670 "Straight Waveguide" sch_x=111 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8336 N$16671 N$16672 "Straight Waveguide" sch_x=111 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8337 N$16673 N$16674 "Straight Waveguide" sch_x=111 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8338 N$16675 N$16676 "Straight Waveguide" sch_x=111 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8339 N$16677 N$16678 "Straight Waveguide" sch_x=111 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8340 N$16679 N$16680 "Straight Waveguide" sch_x=111 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8341 N$16681 N$16682 "Straight Waveguide" sch_x=111 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8342 N$16683 N$16684 "Straight Waveguide" sch_x=111 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8343 N$16685 N$16686 "Straight Waveguide" sch_x=111 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8344 N$16687 N$16688 "Straight Waveguide" sch_x=111 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8345 N$16689 N$16690 "Straight Waveguide" sch_x=109 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8346 N$16691 N$16692 "Straight Waveguide" sch_x=109 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8347 N$16693 N$16694 "Straight Waveguide" sch_x=109 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8348 N$16695 N$16696 "Straight Waveguide" sch_x=109 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8349 N$16697 N$16698 "Straight Waveguide" sch_x=109 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8350 N$16699 N$16700 "Straight Waveguide" sch_x=109 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8351 N$16701 N$16702 "Straight Waveguide" sch_x=109 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8352 N$16703 N$16704 "Straight Waveguide" sch_x=109 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8353 N$16705 N$16706 "Straight Waveguide" sch_x=109 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8354 N$16707 N$16708 "Straight Waveguide" sch_x=109 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8355 N$16709 N$16710 "Straight Waveguide" sch_x=109 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8356 N$16711 N$16712 "Straight Waveguide" sch_x=109 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8357 N$16713 N$16714 "Straight Waveguide" sch_x=109 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8358 N$16715 N$16716 "Straight Waveguide" sch_x=109 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8359 N$16717 N$16718 "Straight Waveguide" sch_x=109 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8360 N$16719 N$16720 "Straight Waveguide" sch_x=109 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8361 N$16721 N$16722 "Straight Waveguide" sch_x=109 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8362 N$16723 N$16724 "Straight Waveguide" sch_x=109 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8363 N$16725 N$16726 "Straight Waveguide" sch_x=109 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8364 N$16727 N$16728 "Straight Waveguide" sch_x=109 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8365 N$16729 N$16730 "Straight Waveguide" sch_x=109 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8366 N$16731 N$16732 "Straight Waveguide" sch_x=109 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8367 N$16733 N$16734 "Straight Waveguide" sch_x=109 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8368 N$16735 N$16736 "Straight Waveguide" sch_x=109 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8369 N$16737 N$16738 "Straight Waveguide" sch_x=109 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8370 N$16739 N$16740 "Straight Waveguide" sch_x=109 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8371 N$16741 N$16742 "Straight Waveguide" sch_x=109 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8372 N$16743 N$16744 "Straight Waveguide" sch_x=109 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8373 N$16745 N$16746 "Straight Waveguide" sch_x=109 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8374 N$16747 N$16748 "Straight Waveguide" sch_x=109 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8375 N$16749 N$16750 "Straight Waveguide" sch_x=109 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8376 N$16751 N$16752 "Straight Waveguide" sch_x=109 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8377 N$16753 N$16754 "Straight Waveguide" sch_x=109 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8378 N$16755 N$16756 "Straight Waveguide" sch_x=109 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8379 N$16757 N$16758 "Straight Waveguide" sch_x=109 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8380 N$16759 N$16760 "Straight Waveguide" sch_x=109 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8381 N$16761 N$16762 "Straight Waveguide" sch_x=109 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8382 N$16763 N$16764 "Straight Waveguide" sch_x=109 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8383 N$16765 N$16766 "Straight Waveguide" sch_x=109 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8384 N$16767 N$16768 "Straight Waveguide" sch_x=109 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8385 N$16769 N$16770 "Straight Waveguide" sch_x=109 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8386 N$16771 N$16772 "Straight Waveguide" sch_x=109 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8387 N$16773 N$16774 "Straight Waveguide" sch_x=109 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8388 N$16775 N$16776 "Straight Waveguide" sch_x=109 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8389 N$16777 N$16778 "Straight Waveguide" sch_x=109 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8390 N$16779 N$16780 "Straight Waveguide" sch_x=109 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8391 N$16781 N$16782 "Straight Waveguide" sch_x=107 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8392 N$16783 N$16784 "Straight Waveguide" sch_x=107 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8393 N$16785 N$16786 "Straight Waveguide" sch_x=107 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8394 N$16787 N$16788 "Straight Waveguide" sch_x=107 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8395 N$16789 N$16790 "Straight Waveguide" sch_x=107 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8396 N$16791 N$16792 "Straight Waveguide" sch_x=107 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8397 N$16793 N$16794 "Straight Waveguide" sch_x=107 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8398 N$16795 N$16796 "Straight Waveguide" sch_x=107 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8399 N$16797 N$16798 "Straight Waveguide" sch_x=107 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8400 N$16799 N$16800 "Straight Waveguide" sch_x=107 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8401 N$16801 N$16802 "Straight Waveguide" sch_x=107 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8402 N$16803 N$16804 "Straight Waveguide" sch_x=107 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8403 N$16805 N$16806 "Straight Waveguide" sch_x=107 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8404 N$16807 N$16808 "Straight Waveguide" sch_x=107 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8405 N$16809 N$16810 "Straight Waveguide" sch_x=107 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8406 N$16811 N$16812 "Straight Waveguide" sch_x=107 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8407 N$16813 N$16814 "Straight Waveguide" sch_x=107 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8408 N$16815 N$16816 "Straight Waveguide" sch_x=107 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8409 N$16817 N$16818 "Straight Waveguide" sch_x=107 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8410 N$16819 N$16820 "Straight Waveguide" sch_x=107 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8411 N$16821 N$16822 "Straight Waveguide" sch_x=107 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8412 N$16823 N$16824 "Straight Waveguide" sch_x=107 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8413 N$16825 N$16826 "Straight Waveguide" sch_x=107 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8414 N$16827 N$16828 "Straight Waveguide" sch_x=107 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8415 N$16829 N$16830 "Straight Waveguide" sch_x=107 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8416 N$16831 N$16832 "Straight Waveguide" sch_x=107 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8417 N$16833 N$16834 "Straight Waveguide" sch_x=107 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8418 N$16835 N$16836 "Straight Waveguide" sch_x=107 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8419 N$16837 N$16838 "Straight Waveguide" sch_x=107 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8420 N$16839 N$16840 "Straight Waveguide" sch_x=107 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8421 N$16841 N$16842 "Straight Waveguide" sch_x=107 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8422 N$16843 N$16844 "Straight Waveguide" sch_x=107 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8423 N$16845 N$16846 "Straight Waveguide" sch_x=107 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8424 N$16847 N$16848 "Straight Waveguide" sch_x=107 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8425 N$16849 N$16850 "Straight Waveguide" sch_x=107 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8426 N$16851 N$16852 "Straight Waveguide" sch_x=107 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8427 N$16853 N$16854 "Straight Waveguide" sch_x=107 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8428 N$16855 N$16856 "Straight Waveguide" sch_x=107 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8429 N$16857 N$16858 "Straight Waveguide" sch_x=107 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8430 N$16859 N$16860 "Straight Waveguide" sch_x=107 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8431 N$16861 N$16862 "Straight Waveguide" sch_x=107 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8432 N$16863 N$16864 "Straight Waveguide" sch_x=107 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8433 N$16865 N$16866 "Straight Waveguide" sch_x=107 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8434 N$16867 N$16868 "Straight Waveguide" sch_x=107 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8435 N$16869 N$16870 "Straight Waveguide" sch_x=105 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8436 N$16871 N$16872 "Straight Waveguide" sch_x=105 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8437 N$16873 N$16874 "Straight Waveguide" sch_x=105 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8438 N$16875 N$16876 "Straight Waveguide" sch_x=105 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8439 N$16877 N$16878 "Straight Waveguide" sch_x=105 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8440 N$16879 N$16880 "Straight Waveguide" sch_x=105 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8441 N$16881 N$16882 "Straight Waveguide" sch_x=105 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8442 N$16883 N$16884 "Straight Waveguide" sch_x=105 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8443 N$16885 N$16886 "Straight Waveguide" sch_x=105 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8444 N$16887 N$16888 "Straight Waveguide" sch_x=105 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8445 N$16889 N$16890 "Straight Waveguide" sch_x=105 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8446 N$16891 N$16892 "Straight Waveguide" sch_x=105 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8447 N$16893 N$16894 "Straight Waveguide" sch_x=105 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8448 N$16895 N$16896 "Straight Waveguide" sch_x=105 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8449 N$16897 N$16898 "Straight Waveguide" sch_x=105 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8450 N$16899 N$16900 "Straight Waveguide" sch_x=105 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8451 N$16901 N$16902 "Straight Waveguide" sch_x=105 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8452 N$16903 N$16904 "Straight Waveguide" sch_x=105 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8453 N$16905 N$16906 "Straight Waveguide" sch_x=105 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8454 N$16907 N$16908 "Straight Waveguide" sch_x=105 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8455 N$16909 N$16910 "Straight Waveguide" sch_x=105 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8456 N$16911 N$16912 "Straight Waveguide" sch_x=105 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8457 N$16913 N$16914 "Straight Waveguide" sch_x=105 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8458 N$16915 N$16916 "Straight Waveguide" sch_x=105 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8459 N$16917 N$16918 "Straight Waveguide" sch_x=105 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8460 N$16919 N$16920 "Straight Waveguide" sch_x=105 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8461 N$16921 N$16922 "Straight Waveguide" sch_x=105 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8462 N$16923 N$16924 "Straight Waveguide" sch_x=105 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8463 N$16925 N$16926 "Straight Waveguide" sch_x=105 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8464 N$16927 N$16928 "Straight Waveguide" sch_x=105 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8465 N$16929 N$16930 "Straight Waveguide" sch_x=105 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8466 N$16931 N$16932 "Straight Waveguide" sch_x=105 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8467 N$16933 N$16934 "Straight Waveguide" sch_x=105 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8468 N$16935 N$16936 "Straight Waveguide" sch_x=105 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8469 N$16937 N$16938 "Straight Waveguide" sch_x=105 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8470 N$16939 N$16940 "Straight Waveguide" sch_x=105 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8471 N$16941 N$16942 "Straight Waveguide" sch_x=105 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8472 N$16943 N$16944 "Straight Waveguide" sch_x=105 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8473 N$16945 N$16946 "Straight Waveguide" sch_x=105 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8474 N$16947 N$16948 "Straight Waveguide" sch_x=105 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8475 N$16949 N$16950 "Straight Waveguide" sch_x=105 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8476 N$16951 N$16952 "Straight Waveguide" sch_x=105 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8477 N$16953 N$16954 "Straight Waveguide" sch_x=103 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8478 N$16955 N$16956 "Straight Waveguide" sch_x=103 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8479 N$16957 N$16958 "Straight Waveguide" sch_x=103 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8480 N$16959 N$16960 "Straight Waveguide" sch_x=103 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8481 N$16961 N$16962 "Straight Waveguide" sch_x=103 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8482 N$16963 N$16964 "Straight Waveguide" sch_x=103 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8483 N$16965 N$16966 "Straight Waveguide" sch_x=103 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8484 N$16967 N$16968 "Straight Waveguide" sch_x=103 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8485 N$16969 N$16970 "Straight Waveguide" sch_x=103 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8486 N$16971 N$16972 "Straight Waveguide" sch_x=103 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8487 N$16973 N$16974 "Straight Waveguide" sch_x=103 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8488 N$16975 N$16976 "Straight Waveguide" sch_x=103 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8489 N$16977 N$16978 "Straight Waveguide" sch_x=103 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8490 N$16979 N$16980 "Straight Waveguide" sch_x=103 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8491 N$16981 N$16982 "Straight Waveguide" sch_x=103 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8492 N$16983 N$16984 "Straight Waveguide" sch_x=103 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8493 N$16985 N$16986 "Straight Waveguide" sch_x=103 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8494 N$16987 N$16988 "Straight Waveguide" sch_x=103 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8495 N$16989 N$16990 "Straight Waveguide" sch_x=103 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8496 N$16991 N$16992 "Straight Waveguide" sch_x=103 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8497 N$16993 N$16994 "Straight Waveguide" sch_x=103 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8498 N$16995 N$16996 "Straight Waveguide" sch_x=103 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8499 N$16997 N$16998 "Straight Waveguide" sch_x=103 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8500 N$16999 N$17000 "Straight Waveguide" sch_x=103 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8501 N$17001 N$17002 "Straight Waveguide" sch_x=103 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8502 N$17003 N$17004 "Straight Waveguide" sch_x=103 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8503 N$17005 N$17006 "Straight Waveguide" sch_x=103 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8504 N$17007 N$17008 "Straight Waveguide" sch_x=103 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8505 N$17009 N$17010 "Straight Waveguide" sch_x=103 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8506 N$17011 N$17012 "Straight Waveguide" sch_x=103 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8507 N$17013 N$17014 "Straight Waveguide" sch_x=103 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8508 N$17015 N$17016 "Straight Waveguide" sch_x=103 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8509 N$17017 N$17018 "Straight Waveguide" sch_x=103 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8510 N$17019 N$17020 "Straight Waveguide" sch_x=103 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8511 N$17021 N$17022 "Straight Waveguide" sch_x=103 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8512 N$17023 N$17024 "Straight Waveguide" sch_x=103 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8513 N$17025 N$17026 "Straight Waveguide" sch_x=103 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8514 N$17027 N$17028 "Straight Waveguide" sch_x=103 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8515 N$17029 N$17030 "Straight Waveguide" sch_x=103 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8516 N$17031 N$17032 "Straight Waveguide" sch_x=103 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8517 N$17033 N$17034 "Straight Waveguide" sch_x=101 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8518 N$17035 N$17036 "Straight Waveguide" sch_x=101 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8519 N$17037 N$17038 "Straight Waveguide" sch_x=101 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8520 N$17039 N$17040 "Straight Waveguide" sch_x=101 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8521 N$17041 N$17042 "Straight Waveguide" sch_x=101 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8522 N$17043 N$17044 "Straight Waveguide" sch_x=101 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8523 N$17045 N$17046 "Straight Waveguide" sch_x=101 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8524 N$17047 N$17048 "Straight Waveguide" sch_x=101 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8525 N$17049 N$17050 "Straight Waveguide" sch_x=101 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8526 N$17051 N$17052 "Straight Waveguide" sch_x=101 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8527 N$17053 N$17054 "Straight Waveguide" sch_x=101 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8528 N$17055 N$17056 "Straight Waveguide" sch_x=101 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8529 N$17057 N$17058 "Straight Waveguide" sch_x=101 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8530 N$17059 N$17060 "Straight Waveguide" sch_x=101 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8531 N$17061 N$17062 "Straight Waveguide" sch_x=101 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8532 N$17063 N$17064 "Straight Waveguide" sch_x=101 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8533 N$17065 N$17066 "Straight Waveguide" sch_x=101 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8534 N$17067 N$17068 "Straight Waveguide" sch_x=101 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8535 N$17069 N$17070 "Straight Waveguide" sch_x=101 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8536 N$17071 N$17072 "Straight Waveguide" sch_x=101 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8537 N$17073 N$17074 "Straight Waveguide" sch_x=101 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8538 N$17075 N$17076 "Straight Waveguide" sch_x=101 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8539 N$17077 N$17078 "Straight Waveguide" sch_x=101 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8540 N$17079 N$17080 "Straight Waveguide" sch_x=101 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8541 N$17081 N$17082 "Straight Waveguide" sch_x=101 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8542 N$17083 N$17084 "Straight Waveguide" sch_x=101 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8543 N$17085 N$17086 "Straight Waveguide" sch_x=101 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8544 N$17087 N$17088 "Straight Waveguide" sch_x=101 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8545 N$17089 N$17090 "Straight Waveguide" sch_x=101 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8546 N$17091 N$17092 "Straight Waveguide" sch_x=101 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8547 N$17093 N$17094 "Straight Waveguide" sch_x=101 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8548 N$17095 N$17096 "Straight Waveguide" sch_x=101 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8549 N$17097 N$17098 "Straight Waveguide" sch_x=101 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8550 N$17099 N$17100 "Straight Waveguide" sch_x=101 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8551 N$17101 N$17102 "Straight Waveguide" sch_x=101 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8552 N$17103 N$17104 "Straight Waveguide" sch_x=101 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8553 N$17105 N$17106 "Straight Waveguide" sch_x=101 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8554 N$17107 N$17108 "Straight Waveguide" sch_x=101 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8555 N$17109 N$17110 "Straight Waveguide" sch_x=99 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8556 N$17111 N$17112 "Straight Waveguide" sch_x=99 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8557 N$17113 N$17114 "Straight Waveguide" sch_x=99 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8558 N$17115 N$17116 "Straight Waveguide" sch_x=99 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8559 N$17117 N$17118 "Straight Waveguide" sch_x=99 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8560 N$17119 N$17120 "Straight Waveguide" sch_x=99 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8561 N$17121 N$17122 "Straight Waveguide" sch_x=99 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8562 N$17123 N$17124 "Straight Waveguide" sch_x=99 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8563 N$17125 N$17126 "Straight Waveguide" sch_x=99 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8564 N$17127 N$17128 "Straight Waveguide" sch_x=99 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8565 N$17129 N$17130 "Straight Waveguide" sch_x=99 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8566 N$17131 N$17132 "Straight Waveguide" sch_x=99 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8567 N$17133 N$17134 "Straight Waveguide" sch_x=99 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8568 N$17135 N$17136 "Straight Waveguide" sch_x=99 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8569 N$17137 N$17138 "Straight Waveguide" sch_x=99 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8570 N$17139 N$17140 "Straight Waveguide" sch_x=99 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8571 N$17141 N$17142 "Straight Waveguide" sch_x=99 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8572 N$17143 N$17144 "Straight Waveguide" sch_x=99 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8573 N$17145 N$17146 "Straight Waveguide" sch_x=99 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8574 N$17147 N$17148 "Straight Waveguide" sch_x=99 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8575 N$17149 N$17150 "Straight Waveguide" sch_x=99 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8576 N$17151 N$17152 "Straight Waveguide" sch_x=99 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8577 N$17153 N$17154 "Straight Waveguide" sch_x=99 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8578 N$17155 N$17156 "Straight Waveguide" sch_x=99 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8579 N$17157 N$17158 "Straight Waveguide" sch_x=99 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8580 N$17159 N$17160 "Straight Waveguide" sch_x=99 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8581 N$17161 N$17162 "Straight Waveguide" sch_x=99 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8582 N$17163 N$17164 "Straight Waveguide" sch_x=99 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8583 N$17165 N$17166 "Straight Waveguide" sch_x=99 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8584 N$17167 N$17168 "Straight Waveguide" sch_x=99 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8585 N$17169 N$17170 "Straight Waveguide" sch_x=99 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8586 N$17171 N$17172 "Straight Waveguide" sch_x=99 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8587 N$17173 N$17174 "Straight Waveguide" sch_x=99 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8588 N$17175 N$17176 "Straight Waveguide" sch_x=99 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8589 N$17177 N$17178 "Straight Waveguide" sch_x=99 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8590 N$17179 N$17180 "Straight Waveguide" sch_x=99 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8591 N$17181 N$17182 "Straight Waveguide" sch_x=97 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8592 N$17183 N$17184 "Straight Waveguide" sch_x=97 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8593 N$17185 N$17186 "Straight Waveguide" sch_x=97 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8594 N$17187 N$17188 "Straight Waveguide" sch_x=97 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8595 N$17189 N$17190 "Straight Waveguide" sch_x=97 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8596 N$17191 N$17192 "Straight Waveguide" sch_x=97 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8597 N$17193 N$17194 "Straight Waveguide" sch_x=97 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8598 N$17195 N$17196 "Straight Waveguide" sch_x=97 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8599 N$17197 N$17198 "Straight Waveguide" sch_x=97 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8600 N$17199 N$17200 "Straight Waveguide" sch_x=97 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8601 N$17201 N$17202 "Straight Waveguide" sch_x=97 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8602 N$17203 N$17204 "Straight Waveguide" sch_x=97 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8603 N$17205 N$17206 "Straight Waveguide" sch_x=97 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8604 N$17207 N$17208 "Straight Waveguide" sch_x=97 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8605 N$17209 N$17210 "Straight Waveguide" sch_x=97 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8606 N$17211 N$17212 "Straight Waveguide" sch_x=97 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8607 N$17213 N$17214 "Straight Waveguide" sch_x=97 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8608 N$17215 N$17216 "Straight Waveguide" sch_x=97 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8609 N$17217 N$17218 "Straight Waveguide" sch_x=97 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8610 N$17219 N$17220 "Straight Waveguide" sch_x=97 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8611 N$17221 N$17222 "Straight Waveguide" sch_x=97 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8612 N$17223 N$17224 "Straight Waveguide" sch_x=97 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8613 N$17225 N$17226 "Straight Waveguide" sch_x=97 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8614 N$17227 N$17228 "Straight Waveguide" sch_x=97 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8615 N$17229 N$17230 "Straight Waveguide" sch_x=97 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8616 N$17231 N$17232 "Straight Waveguide" sch_x=97 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8617 N$17233 N$17234 "Straight Waveguide" sch_x=97 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8618 N$17235 N$17236 "Straight Waveguide" sch_x=97 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8619 N$17237 N$17238 "Straight Waveguide" sch_x=97 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8620 N$17239 N$17240 "Straight Waveguide" sch_x=97 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8621 N$17241 N$17242 "Straight Waveguide" sch_x=97 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8622 N$17243 N$17244 "Straight Waveguide" sch_x=97 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8623 N$17245 N$17246 "Straight Waveguide" sch_x=97 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8624 N$17247 N$17248 "Straight Waveguide" sch_x=97 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8625 N$17249 N$17250 "Straight Waveguide" sch_x=95 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8626 N$17251 N$17252 "Straight Waveguide" sch_x=95 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8627 N$17253 N$17254 "Straight Waveguide" sch_x=95 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8628 N$17255 N$17256 "Straight Waveguide" sch_x=95 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8629 N$17257 N$17258 "Straight Waveguide" sch_x=95 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8630 N$17259 N$17260 "Straight Waveguide" sch_x=95 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8631 N$17261 N$17262 "Straight Waveguide" sch_x=95 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8632 N$17263 N$17264 "Straight Waveguide" sch_x=95 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8633 N$17265 N$17266 "Straight Waveguide" sch_x=95 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8634 N$17267 N$17268 "Straight Waveguide" sch_x=95 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8635 N$17269 N$17270 "Straight Waveguide" sch_x=95 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8636 N$17271 N$17272 "Straight Waveguide" sch_x=95 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8637 N$17273 N$17274 "Straight Waveguide" sch_x=95 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8638 N$17275 N$17276 "Straight Waveguide" sch_x=95 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8639 N$17277 N$17278 "Straight Waveguide" sch_x=95 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8640 N$17279 N$17280 "Straight Waveguide" sch_x=95 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8641 N$17281 N$17282 "Straight Waveguide" sch_x=95 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8642 N$17283 N$17284 "Straight Waveguide" sch_x=95 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8643 N$17285 N$17286 "Straight Waveguide" sch_x=95 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8644 N$17287 N$17288 "Straight Waveguide" sch_x=95 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8645 N$17289 N$17290 "Straight Waveguide" sch_x=95 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8646 N$17291 N$17292 "Straight Waveguide" sch_x=95 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8647 N$17293 N$17294 "Straight Waveguide" sch_x=95 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8648 N$17295 N$17296 "Straight Waveguide" sch_x=95 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8649 N$17297 N$17298 "Straight Waveguide" sch_x=95 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8650 N$17299 N$17300 "Straight Waveguide" sch_x=95 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8651 N$17301 N$17302 "Straight Waveguide" sch_x=95 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8652 N$17303 N$17304 "Straight Waveguide" sch_x=95 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8653 N$17305 N$17306 "Straight Waveguide" sch_x=95 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8654 N$17307 N$17308 "Straight Waveguide" sch_x=95 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8655 N$17309 N$17310 "Straight Waveguide" sch_x=95 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8656 N$17311 N$17312 "Straight Waveguide" sch_x=95 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8657 N$17313 N$17314 "Straight Waveguide" sch_x=93 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8658 N$17315 N$17316 "Straight Waveguide" sch_x=93 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8659 N$17317 N$17318 "Straight Waveguide" sch_x=93 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8660 N$17319 N$17320 "Straight Waveguide" sch_x=93 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8661 N$17321 N$17322 "Straight Waveguide" sch_x=93 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8662 N$17323 N$17324 "Straight Waveguide" sch_x=93 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8663 N$17325 N$17326 "Straight Waveguide" sch_x=93 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8664 N$17327 N$17328 "Straight Waveguide" sch_x=93 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8665 N$17329 N$17330 "Straight Waveguide" sch_x=93 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8666 N$17331 N$17332 "Straight Waveguide" sch_x=93 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8667 N$17333 N$17334 "Straight Waveguide" sch_x=93 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8668 N$17335 N$17336 "Straight Waveguide" sch_x=93 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8669 N$17337 N$17338 "Straight Waveguide" sch_x=93 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8670 N$17339 N$17340 "Straight Waveguide" sch_x=93 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8671 N$17341 N$17342 "Straight Waveguide" sch_x=93 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8672 N$17343 N$17344 "Straight Waveguide" sch_x=93 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8673 N$17345 N$17346 "Straight Waveguide" sch_x=93 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8674 N$17347 N$17348 "Straight Waveguide" sch_x=93 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8675 N$17349 N$17350 "Straight Waveguide" sch_x=93 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8676 N$17351 N$17352 "Straight Waveguide" sch_x=93 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8677 N$17353 N$17354 "Straight Waveguide" sch_x=93 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8678 N$17355 N$17356 "Straight Waveguide" sch_x=93 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8679 N$17357 N$17358 "Straight Waveguide" sch_x=93 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8680 N$17359 N$17360 "Straight Waveguide" sch_x=93 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8681 N$17361 N$17362 "Straight Waveguide" sch_x=93 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8682 N$17363 N$17364 "Straight Waveguide" sch_x=93 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8683 N$17365 N$17366 "Straight Waveguide" sch_x=93 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8684 N$17367 N$17368 "Straight Waveguide" sch_x=93 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8685 N$17369 N$17370 "Straight Waveguide" sch_x=93 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8686 N$17371 N$17372 "Straight Waveguide" sch_x=93 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8687 N$17373 N$17374 "Straight Waveguide" sch_x=91 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8688 N$17375 N$17376 "Straight Waveguide" sch_x=91 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8689 N$17377 N$17378 "Straight Waveguide" sch_x=91 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8690 N$17379 N$17380 "Straight Waveguide" sch_x=91 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8691 N$17381 N$17382 "Straight Waveguide" sch_x=91 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8692 N$17383 N$17384 "Straight Waveguide" sch_x=91 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8693 N$17385 N$17386 "Straight Waveguide" sch_x=91 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8694 N$17387 N$17388 "Straight Waveguide" sch_x=91 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8695 N$17389 N$17390 "Straight Waveguide" sch_x=91 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8696 N$17391 N$17392 "Straight Waveguide" sch_x=91 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8697 N$17393 N$17394 "Straight Waveguide" sch_x=91 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8698 N$17395 N$17396 "Straight Waveguide" sch_x=91 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8699 N$17397 N$17398 "Straight Waveguide" sch_x=91 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8700 N$17399 N$17400 "Straight Waveguide" sch_x=91 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8701 N$17401 N$17402 "Straight Waveguide" sch_x=91 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8702 N$17403 N$17404 "Straight Waveguide" sch_x=91 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8703 N$17405 N$17406 "Straight Waveguide" sch_x=91 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8704 N$17407 N$17408 "Straight Waveguide" sch_x=91 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8705 N$17409 N$17410 "Straight Waveguide" sch_x=91 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8706 N$17411 N$17412 "Straight Waveguide" sch_x=91 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8707 N$17413 N$17414 "Straight Waveguide" sch_x=91 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8708 N$17415 N$17416 "Straight Waveguide" sch_x=91 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8709 N$17417 N$17418 "Straight Waveguide" sch_x=91 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8710 N$17419 N$17420 "Straight Waveguide" sch_x=91 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8711 N$17421 N$17422 "Straight Waveguide" sch_x=91 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8712 N$17423 N$17424 "Straight Waveguide" sch_x=91 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8713 N$17425 N$17426 "Straight Waveguide" sch_x=91 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8714 N$17427 N$17428 "Straight Waveguide" sch_x=91 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8715 N$17429 N$17430 "Straight Waveguide" sch_x=89 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8716 N$17431 N$17432 "Straight Waveguide" sch_x=89 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8717 N$17433 N$17434 "Straight Waveguide" sch_x=89 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8718 N$17435 N$17436 "Straight Waveguide" sch_x=89 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8719 N$17437 N$17438 "Straight Waveguide" sch_x=89 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8720 N$17439 N$17440 "Straight Waveguide" sch_x=89 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8721 N$17441 N$17442 "Straight Waveguide" sch_x=89 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8722 N$17443 N$17444 "Straight Waveguide" sch_x=89 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8723 N$17445 N$17446 "Straight Waveguide" sch_x=89 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8724 N$17447 N$17448 "Straight Waveguide" sch_x=89 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8725 N$17449 N$17450 "Straight Waveguide" sch_x=89 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8726 N$17451 N$17452 "Straight Waveguide" sch_x=89 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8727 N$17453 N$17454 "Straight Waveguide" sch_x=89 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8728 N$17455 N$17456 "Straight Waveguide" sch_x=89 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8729 N$17457 N$17458 "Straight Waveguide" sch_x=89 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8730 N$17459 N$17460 "Straight Waveguide" sch_x=89 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8731 N$17461 N$17462 "Straight Waveguide" sch_x=89 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8732 N$17463 N$17464 "Straight Waveguide" sch_x=89 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8733 N$17465 N$17466 "Straight Waveguide" sch_x=89 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8734 N$17467 N$17468 "Straight Waveguide" sch_x=89 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8735 N$17469 N$17470 "Straight Waveguide" sch_x=89 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8736 N$17471 N$17472 "Straight Waveguide" sch_x=89 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8737 N$17473 N$17474 "Straight Waveguide" sch_x=89 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8738 N$17475 N$17476 "Straight Waveguide" sch_x=89 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8739 N$17477 N$17478 "Straight Waveguide" sch_x=89 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8740 N$17479 N$17480 "Straight Waveguide" sch_x=89 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8741 N$17481 N$17482 "Straight Waveguide" sch_x=87 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8742 N$17483 N$17484 "Straight Waveguide" sch_x=87 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8743 N$17485 N$17486 "Straight Waveguide" sch_x=87 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8744 N$17487 N$17488 "Straight Waveguide" sch_x=87 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8745 N$17489 N$17490 "Straight Waveguide" sch_x=87 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8746 N$17491 N$17492 "Straight Waveguide" sch_x=87 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8747 N$17493 N$17494 "Straight Waveguide" sch_x=87 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8748 N$17495 N$17496 "Straight Waveguide" sch_x=87 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8749 N$17497 N$17498 "Straight Waveguide" sch_x=87 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8750 N$17499 N$17500 "Straight Waveguide" sch_x=87 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8751 N$17501 N$17502 "Straight Waveguide" sch_x=87 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8752 N$17503 N$17504 "Straight Waveguide" sch_x=87 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8753 N$17505 N$17506 "Straight Waveguide" sch_x=87 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8754 N$17507 N$17508 "Straight Waveguide" sch_x=87 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8755 N$17509 N$17510 "Straight Waveguide" sch_x=87 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8756 N$17511 N$17512 "Straight Waveguide" sch_x=87 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8757 N$17513 N$17514 "Straight Waveguide" sch_x=87 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8758 N$17515 N$17516 "Straight Waveguide" sch_x=87 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8759 N$17517 N$17518 "Straight Waveguide" sch_x=87 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8760 N$17519 N$17520 "Straight Waveguide" sch_x=87 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8761 N$17521 N$17522 "Straight Waveguide" sch_x=87 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8762 N$17523 N$17524 "Straight Waveguide" sch_x=87 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8763 N$17525 N$17526 "Straight Waveguide" sch_x=87 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8764 N$17527 N$17528 "Straight Waveguide" sch_x=87 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8765 N$17529 N$17530 "Straight Waveguide" sch_x=85 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8766 N$17531 N$17532 "Straight Waveguide" sch_x=85 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8767 N$17533 N$17534 "Straight Waveguide" sch_x=85 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8768 N$17535 N$17536 "Straight Waveguide" sch_x=85 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8769 N$17537 N$17538 "Straight Waveguide" sch_x=85 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8770 N$17539 N$17540 "Straight Waveguide" sch_x=85 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8771 N$17541 N$17542 "Straight Waveguide" sch_x=85 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8772 N$17543 N$17544 "Straight Waveguide" sch_x=85 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8773 N$17545 N$17546 "Straight Waveguide" sch_x=85 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8774 N$17547 N$17548 "Straight Waveguide" sch_x=85 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8775 N$17549 N$17550 "Straight Waveguide" sch_x=85 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8776 N$17551 N$17552 "Straight Waveguide" sch_x=85 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8777 N$17553 N$17554 "Straight Waveguide" sch_x=85 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8778 N$17555 N$17556 "Straight Waveguide" sch_x=85 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8779 N$17557 N$17558 "Straight Waveguide" sch_x=85 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8780 N$17559 N$17560 "Straight Waveguide" sch_x=85 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8781 N$17561 N$17562 "Straight Waveguide" sch_x=85 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8782 N$17563 N$17564 "Straight Waveguide" sch_x=85 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8783 N$17565 N$17566 "Straight Waveguide" sch_x=85 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8784 N$17567 N$17568 "Straight Waveguide" sch_x=85 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8785 N$17569 N$17570 "Straight Waveguide" sch_x=85 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8786 N$17571 N$17572 "Straight Waveguide" sch_x=85 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8787 N$17573 N$17574 "Straight Waveguide" sch_x=83 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8788 N$17575 N$17576 "Straight Waveguide" sch_x=83 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8789 N$17577 N$17578 "Straight Waveguide" sch_x=83 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8790 N$17579 N$17580 "Straight Waveguide" sch_x=83 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8791 N$17581 N$17582 "Straight Waveguide" sch_x=83 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8792 N$17583 N$17584 "Straight Waveguide" sch_x=83 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8793 N$17585 N$17586 "Straight Waveguide" sch_x=83 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8794 N$17587 N$17588 "Straight Waveguide" sch_x=83 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8795 N$17589 N$17590 "Straight Waveguide" sch_x=83 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8796 N$17591 N$17592 "Straight Waveguide" sch_x=83 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8797 N$17593 N$17594 "Straight Waveguide" sch_x=83 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8798 N$17595 N$17596 "Straight Waveguide" sch_x=83 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8799 N$17597 N$17598 "Straight Waveguide" sch_x=83 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8800 N$17599 N$17600 "Straight Waveguide" sch_x=83 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8801 N$17601 N$17602 "Straight Waveguide" sch_x=83 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8802 N$17603 N$17604 "Straight Waveguide" sch_x=83 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8803 N$17605 N$17606 "Straight Waveguide" sch_x=83 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8804 N$17607 N$17608 "Straight Waveguide" sch_x=83 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8805 N$17609 N$17610 "Straight Waveguide" sch_x=83 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8806 N$17611 N$17612 "Straight Waveguide" sch_x=83 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8807 N$17613 N$17614 "Straight Waveguide" sch_x=81 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8808 N$17615 N$17616 "Straight Waveguide" sch_x=81 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8809 N$17617 N$17618 "Straight Waveguide" sch_x=81 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8810 N$17619 N$17620 "Straight Waveguide" sch_x=81 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8811 N$17621 N$17622 "Straight Waveguide" sch_x=81 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8812 N$17623 N$17624 "Straight Waveguide" sch_x=81 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8813 N$17625 N$17626 "Straight Waveguide" sch_x=81 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8814 N$17627 N$17628 "Straight Waveguide" sch_x=81 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8815 N$17629 N$17630 "Straight Waveguide" sch_x=81 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8816 N$17631 N$17632 "Straight Waveguide" sch_x=81 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8817 N$17633 N$17634 "Straight Waveguide" sch_x=81 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8818 N$17635 N$17636 "Straight Waveguide" sch_x=81 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8819 N$17637 N$17638 "Straight Waveguide" sch_x=81 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8820 N$17639 N$17640 "Straight Waveguide" sch_x=81 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8821 N$17641 N$17642 "Straight Waveguide" sch_x=81 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8822 N$17643 N$17644 "Straight Waveguide" sch_x=81 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8823 N$17645 N$17646 "Straight Waveguide" sch_x=81 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8824 N$17647 N$17648 "Straight Waveguide" sch_x=81 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8825 N$17649 N$17650 "Straight Waveguide" sch_x=79 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8826 N$17651 N$17652 "Straight Waveguide" sch_x=79 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8827 N$17653 N$17654 "Straight Waveguide" sch_x=79 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8828 N$17655 N$17656 "Straight Waveguide" sch_x=79 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8829 N$17657 N$17658 "Straight Waveguide" sch_x=79 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8830 N$17659 N$17660 "Straight Waveguide" sch_x=79 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8831 N$17661 N$17662 "Straight Waveguide" sch_x=79 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8832 N$17663 N$17664 "Straight Waveguide" sch_x=79 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8833 N$17665 N$17666 "Straight Waveguide" sch_x=79 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8834 N$17667 N$17668 "Straight Waveguide" sch_x=79 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8835 N$17669 N$17670 "Straight Waveguide" sch_x=79 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8836 N$17671 N$17672 "Straight Waveguide" sch_x=79 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8837 N$17673 N$17674 "Straight Waveguide" sch_x=79 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8838 N$17675 N$17676 "Straight Waveguide" sch_x=79 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8839 N$17677 N$17678 "Straight Waveguide" sch_x=79 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8840 N$17679 N$17680 "Straight Waveguide" sch_x=79 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8841 N$17681 N$17682 "Straight Waveguide" sch_x=77 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8842 N$17683 N$17684 "Straight Waveguide" sch_x=77 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8843 N$17685 N$17686 "Straight Waveguide" sch_x=77 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8844 N$17687 N$17688 "Straight Waveguide" sch_x=77 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8845 N$17689 N$17690 "Straight Waveguide" sch_x=77 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8846 N$17691 N$17692 "Straight Waveguide" sch_x=77 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8847 N$17693 N$17694 "Straight Waveguide" sch_x=77 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8848 N$17695 N$17696 "Straight Waveguide" sch_x=77 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8849 N$17697 N$17698 "Straight Waveguide" sch_x=77 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8850 N$17699 N$17700 "Straight Waveguide" sch_x=77 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8851 N$17701 N$17702 "Straight Waveguide" sch_x=77 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8852 N$17703 N$17704 "Straight Waveguide" sch_x=77 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8853 N$17705 N$17706 "Straight Waveguide" sch_x=77 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8854 N$17707 N$17708 "Straight Waveguide" sch_x=77 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8855 N$17709 N$17710 "Straight Waveguide" sch_x=75 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8856 N$17711 N$17712 "Straight Waveguide" sch_x=75 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8857 N$17713 N$17714 "Straight Waveguide" sch_x=75 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8858 N$17715 N$17716 "Straight Waveguide" sch_x=75 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8859 N$17717 N$17718 "Straight Waveguide" sch_x=75 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8860 N$17719 N$17720 "Straight Waveguide" sch_x=75 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8861 N$17721 N$17722 "Straight Waveguide" sch_x=75 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8862 N$17723 N$17724 "Straight Waveguide" sch_x=75 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8863 N$17725 N$17726 "Straight Waveguide" sch_x=75 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8864 N$17727 N$17728 "Straight Waveguide" sch_x=75 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8865 N$17729 N$17730 "Straight Waveguide" sch_x=75 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8866 N$17731 N$17732 "Straight Waveguide" sch_x=75 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8867 N$17733 N$17734 "Straight Waveguide" sch_x=73 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8868 N$17735 N$17736 "Straight Waveguide" sch_x=73 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8869 N$17737 N$17738 "Straight Waveguide" sch_x=73 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8870 N$17739 N$17740 "Straight Waveguide" sch_x=73 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8871 N$17741 N$17742 "Straight Waveguide" sch_x=73 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8872 N$17743 N$17744 "Straight Waveguide" sch_x=73 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8873 N$17745 N$17746 "Straight Waveguide" sch_x=73 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8874 N$17747 N$17748 "Straight Waveguide" sch_x=73 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8875 N$17749 N$17750 "Straight Waveguide" sch_x=73 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8876 N$17751 N$17752 "Straight Waveguide" sch_x=73 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8877 N$17753 N$17754 "Straight Waveguide" sch_x=71 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8878 N$17755 N$17756 "Straight Waveguide" sch_x=71 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8879 N$17757 N$17758 "Straight Waveguide" sch_x=71 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8880 N$17759 N$17760 "Straight Waveguide" sch_x=71 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8881 N$17761 N$17762 "Straight Waveguide" sch_x=71 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8882 N$17763 N$17764 "Straight Waveguide" sch_x=71 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8883 N$17765 N$17766 "Straight Waveguide" sch_x=71 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8884 N$17767 N$17768 "Straight Waveguide" sch_x=71 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8885 N$17769 N$17770 "Straight Waveguide" sch_x=69 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8886 N$17771 N$17772 "Straight Waveguide" sch_x=69 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8887 N$17773 N$17774 "Straight Waveguide" sch_x=69 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8888 N$17775 N$17776 "Straight Waveguide" sch_x=69 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8889 N$17777 N$17778 "Straight Waveguide" sch_x=69 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8890 N$17779 N$17780 "Straight Waveguide" sch_x=69 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8891 N$17781 N$17782 "Straight Waveguide" sch_x=67 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8892 N$17783 N$17784 "Straight Waveguide" sch_x=67 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8893 N$17785 N$17786 "Straight Waveguide" sch_x=67 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8894 N$17787 N$17788 "Straight Waveguide" sch_x=67 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8895 N$17789 N$17790 "Straight Waveguide" sch_x=65 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8896 N$17791 N$17792 "Straight Waveguide" sch_x=65 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8897 N$17794 N$17793 "Straight Waveguide" sch_x=93 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8898 N$17796 N$17795 "Straight Waveguide" sch_x=92 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8899 N$17798 N$17797 "Straight Waveguide" sch_x=91 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8900 N$17800 N$17799 "Straight Waveguide" sch_x=90 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8901 N$17802 N$17801 "Straight Waveguide" sch_x=89 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8902 N$17804 N$17803 "Straight Waveguide" sch_x=88 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8903 N$17806 N$17805 "Straight Waveguide" sch_x=87 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8904 N$17808 N$17807 "Straight Waveguide" sch_x=86 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8905 N$17810 N$17809 "Straight Waveguide" sch_x=85 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8906 N$17812 N$17811 "Straight Waveguide" sch_x=84 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8907 N$17814 N$17813 "Straight Waveguide" sch_x=83 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8908 N$17816 N$17815 "Straight Waveguide" sch_x=82 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8909 N$17818 N$17817 "Straight Waveguide" sch_x=81 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8910 N$17820 N$17819 "Straight Waveguide" sch_x=80 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8911 N$17822 N$17821 "Straight Waveguide" sch_x=79 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8912 N$17824 N$17823 "Straight Waveguide" sch_x=78 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8913 N$17826 N$17825 "Straight Waveguide" sch_x=77 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8914 N$17828 N$17827 "Straight Waveguide" sch_x=76 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8915 N$17830 N$17829 "Straight Waveguide" sch_x=75 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8916 N$17832 N$17831 "Straight Waveguide" sch_x=74 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8917 N$17834 N$17833 "Straight Waveguide" sch_x=73 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8918 N$17836 N$17835 "Straight Waveguide" sch_x=72 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8919 N$17838 N$17837 "Straight Waveguide" sch_x=71 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8920 N$17840 N$17839 "Straight Waveguide" sch_x=70 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8921 N$17842 N$17841 "Straight Waveguide" sch_x=69 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8922 N$17844 N$17843 "Straight Waveguide" sch_x=68 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8923 N$17846 N$17845 "Straight Waveguide" sch_x=67 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8924 N$17848 N$17847 "Straight Waveguide" sch_x=66 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8925 N$17850 N$17849 "Straight Waveguide" sch_x=65 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8926 N$17852 N$17851 "Straight Waveguide" sch_x=64 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8927 N$17854 N$17853 "Straight Waveguide" sch_x=63 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8928 N$17856 N$17855 "Straight Waveguide" sch_x=63 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8929 N$17858 N$17857 "Straight Waveguide" sch_x=64 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8930 N$17860 N$17859 "Straight Waveguide" sch_x=65 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8931 N$17862 N$17861 "Straight Waveguide" sch_x=66 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8932 N$17864 N$17863 "Straight Waveguide" sch_x=67 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8933 N$17866 N$17865 "Straight Waveguide" sch_x=68 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8934 N$17868 N$17867 "Straight Waveguide" sch_x=69 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8935 N$17870 N$17869 "Straight Waveguide" sch_x=70 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8936 N$17872 N$17871 "Straight Waveguide" sch_x=71 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8937 N$17874 N$17873 "Straight Waveguide" sch_x=72 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8938 N$17876 N$17875 "Straight Waveguide" sch_x=73 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8939 N$17878 N$17877 "Straight Waveguide" sch_x=74 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8940 N$17880 N$17879 "Straight Waveguide" sch_x=75 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8941 N$17882 N$17881 "Straight Waveguide" sch_x=76 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8942 N$17884 N$17883 "Straight Waveguide" sch_x=77 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8943 N$17886 N$17885 "Straight Waveguide" sch_x=78 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8944 N$17888 N$17887 "Straight Waveguide" sch_x=79 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8945 N$17890 N$17889 "Straight Waveguide" sch_x=80 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8946 N$17892 N$17891 "Straight Waveguide" sch_x=81 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8947 N$17894 N$17893 "Straight Waveguide" sch_x=82 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8948 N$17896 N$17895 "Straight Waveguide" sch_x=83 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8949 N$17898 N$17897 "Straight Waveguide" sch_x=84 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8950 N$17900 N$17899 "Straight Waveguide" sch_x=85 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8951 N$17902 N$17901 "Straight Waveguide" sch_x=86 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8952 N$17904 N$17903 "Straight Waveguide" sch_x=87 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8953 N$17906 N$17905 "Straight Waveguide" sch_x=88 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8954 N$17908 N$17907 "Straight Waveguide" sch_x=89 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8955 N$17910 N$17909 "Straight Waveguide" sch_x=90 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8956 N$17912 N$17911 "Straight Waveguide" sch_x=91 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8957 N$17914 N$17913 "Straight Waveguide" sch_x=92 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8958 N$17916 N$17915 "Straight Waveguide" sch_x=93 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8959 N$17918 N$17917 "Straight Waveguide" sch_x=94 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8960 N$17920 N$17919 "Straight Waveguide" sch_x=94 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8961 N$17922 N$17921 "Straight Waveguide" sch_x=-253 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8962 N$17924 N$17923 "Straight Waveguide" sch_x=-253 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8963 N$17926 N$17925 "Straight Waveguide" sch_x=-253 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8964 N$17928 N$17927 "Straight Waveguide" sch_x=-253 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8965 N$17930 N$17929 "Straight Waveguide" sch_x=-253 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8966 N$17932 N$17931 "Straight Waveguide" sch_x=-253 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8967 N$17934 N$17933 "Straight Waveguide" sch_x=-253 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8968 N$17936 N$17935 "Straight Waveguide" sch_x=-253 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8969 N$17938 N$17937 "Straight Waveguide" sch_x=-253 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8970 N$17940 N$17939 "Straight Waveguide" sch_x=-253 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8971 N$17942 N$17941 "Straight Waveguide" sch_x=-253 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8972 N$17944 N$17943 "Straight Waveguide" sch_x=-253 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8973 N$17946 N$17945 "Straight Waveguide" sch_x=-253 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8974 N$17948 N$17947 "Straight Waveguide" sch_x=-253 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8975 N$17950 N$17949 "Straight Waveguide" sch_x=-253 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8976 N$17952 N$17951 "Straight Waveguide" sch_x=-253 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8977 N$17954 N$17953 "Straight Waveguide" sch_x=-253 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8978 N$17956 N$17955 "Straight Waveguide" sch_x=-253 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8979 N$17958 N$17957 "Straight Waveguide" sch_x=-253 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8980 N$17960 N$17959 "Straight Waveguide" sch_x=-253 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8981 N$17962 N$17961 "Straight Waveguide" sch_x=-253 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8982 N$17964 N$17963 "Straight Waveguide" sch_x=-253 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8983 N$17966 N$17965 "Straight Waveguide" sch_x=-253 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8984 N$17968 N$17967 "Straight Waveguide" sch_x=-253 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8985 N$17970 N$17969 "Straight Waveguide" sch_x=-253 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8986 N$17972 N$17971 "Straight Waveguide" sch_x=-253 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8987 N$17974 N$17973 "Straight Waveguide" sch_x=-253 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8988 N$17976 N$17975 "Straight Waveguide" sch_x=-253 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8989 N$17978 N$17977 "Straight Waveguide" sch_x=-253 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8990 N$17980 N$17979 "Straight Waveguide" sch_x=-253 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8991 N$17982 N$17981 "Straight Waveguide" sch_x=-253 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8992 N$17984 N$17983 "Straight Waveguide" sch_x=-253 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8993 N$17986 N$17985 "Straight Waveguide" sch_x=-253 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8994 N$17988 N$17987 "Straight Waveguide" sch_x=-253 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8995 N$17990 N$17989 "Straight Waveguide" sch_x=-253 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8996 N$17992 N$17991 "Straight Waveguide" sch_x=-253 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8997 N$17994 N$17993 "Straight Waveguide" sch_x=-253 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8998 N$17996 N$17995 "Straight Waveguide" sch_x=-253 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8999 N$17998 N$17997 "Straight Waveguide" sch_x=-253 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9000 N$18000 N$17999 "Straight Waveguide" sch_x=-253 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9001 N$18002 N$18001 "Straight Waveguide" sch_x=-253 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9002 N$18004 N$18003 "Straight Waveguide" sch_x=-253 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9003 N$18006 N$18005 "Straight Waveguide" sch_x=-253 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9004 N$18008 N$18007 "Straight Waveguide" sch_x=-253 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9005 N$18010 N$18009 "Straight Waveguide" sch_x=-253 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9006 N$18012 N$18011 "Straight Waveguide" sch_x=-253 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9007 N$18014 N$18013 "Straight Waveguide" sch_x=-253 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9008 N$18016 N$18015 "Straight Waveguide" sch_x=-253 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9009 N$18018 N$18017 "Straight Waveguide" sch_x=-253 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9010 N$18020 N$18019 "Straight Waveguide" sch_x=-253 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9011 N$18022 N$18021 "Straight Waveguide" sch_x=-253 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9012 N$18024 N$18023 "Straight Waveguide" sch_x=-253 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9013 N$18026 N$18025 "Straight Waveguide" sch_x=-253 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9014 N$18028 N$18027 "Straight Waveguide" sch_x=-253 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9015 N$18030 N$18029 "Straight Waveguide" sch_x=-253 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9016 N$18032 N$18031 "Straight Waveguide" sch_x=-253 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9017 N$18034 N$18033 "Straight Waveguide" sch_x=-253 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9018 N$18036 N$18035 "Straight Waveguide" sch_x=-253 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9019 N$18038 N$18037 "Straight Waveguide" sch_x=-253 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9020 N$18040 N$18039 "Straight Waveguide" sch_x=-253 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9021 N$18042 N$18041 "Straight Waveguide" sch_x=-253 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9022 N$18044 N$18043 "Straight Waveguide" sch_x=-253 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9023 N$18046 N$18045 "Straight Waveguide" sch_x=-253 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9024 N$18048 N$18047 "Straight Waveguide" sch_x=-253 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9025 N$18050 N$18049 "Straight Waveguide" sch_x=-253 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9026 N$18052 N$18051 "Straight Waveguide" sch_x=-253 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9027 N$18054 N$18053 "Straight Waveguide" sch_x=-253 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9028 N$18056 N$18055 "Straight Waveguide" sch_x=-253 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9029 N$18058 N$18057 "Straight Waveguide" sch_x=-253 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9030 N$18060 N$18059 "Straight Waveguide" sch_x=-253 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9031 N$18062 N$18061 "Straight Waveguide" sch_x=-253 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9032 N$18064 N$18063 "Straight Waveguide" sch_x=-253 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9033 N$18066 N$18065 "Straight Waveguide" sch_x=-253 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9034 N$18068 N$18067 "Straight Waveguide" sch_x=-253 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9035 N$18070 N$18069 "Straight Waveguide" sch_x=-253 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9036 N$18072 N$18071 "Straight Waveguide" sch_x=-253 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9037 N$18074 N$18073 "Straight Waveguide" sch_x=-253 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9038 N$18076 N$18075 "Straight Waveguide" sch_x=-253 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9039 N$18078 N$18077 "Straight Waveguide" sch_x=-253 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9040 N$18080 N$18079 "Straight Waveguide" sch_x=-253 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9041 N$18082 N$18081 "Straight Waveguide" sch_x=-253 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9042 N$18084 N$18083 "Straight Waveguide" sch_x=-253 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9043 N$18086 N$18085 "Straight Waveguide" sch_x=-253 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9044 N$18088 N$18087 "Straight Waveguide" sch_x=-253 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9045 N$18090 N$18089 "Straight Waveguide" sch_x=-253 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9046 N$18092 N$18091 "Straight Waveguide" sch_x=-253 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9047 N$18094 N$18093 "Straight Waveguide" sch_x=-253 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9048 N$18096 N$18095 "Straight Waveguide" sch_x=-253 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9049 N$18098 N$18097 "Straight Waveguide" sch_x=-253 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9050 N$18100 N$18099 "Straight Waveguide" sch_x=-253 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9051 N$18102 N$18101 "Straight Waveguide" sch_x=-253 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9052 N$18104 N$18103 "Straight Waveguide" sch_x=-253 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9053 N$18106 N$18105 "Straight Waveguide" sch_x=-253 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9054 N$18108 N$18107 "Straight Waveguide" sch_x=-253 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9055 N$18110 N$18109 "Straight Waveguide" sch_x=-253 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9056 N$18112 N$18111 "Straight Waveguide" sch_x=-253 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9057 N$18114 N$18113 "Straight Waveguide" sch_x=-253 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9058 N$18116 N$18115 "Straight Waveguide" sch_x=-253 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9059 N$18118 N$18117 "Straight Waveguide" sch_x=-253 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9060 N$18120 N$18119 "Straight Waveguide" sch_x=-253 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9061 N$18122 N$18121 "Straight Waveguide" sch_x=-253 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9062 N$18124 N$18123 "Straight Waveguide" sch_x=-253 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9063 N$18126 N$18125 "Straight Waveguide" sch_x=-253 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9064 N$18128 N$18127 "Straight Waveguide" sch_x=-253 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9065 N$18130 N$18129 "Straight Waveguide" sch_x=-253 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9066 N$18132 N$18131 "Straight Waveguide" sch_x=-253 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9067 N$18134 N$18133 "Straight Waveguide" sch_x=-253 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9068 N$18136 N$18135 "Straight Waveguide" sch_x=-253 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9069 N$18138 N$18137 "Straight Waveguide" sch_x=-253 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9070 N$18140 N$18139 "Straight Waveguide" sch_x=-253 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9071 N$18142 N$18141 "Straight Waveguide" sch_x=-253 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9072 N$18144 N$18143 "Straight Waveguide" sch_x=-253 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9073 N$18146 N$18145 "Straight Waveguide" sch_x=-253 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9074 N$18148 N$18147 "Straight Waveguide" sch_x=-253 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9075 N$18150 N$18149 "Straight Waveguide" sch_x=-253 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9076 N$18152 N$18151 "Straight Waveguide" sch_x=-253 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9077 N$18154 N$18153 "Straight Waveguide" sch_x=-253 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9078 N$18156 N$18155 "Straight Waveguide" sch_x=-253 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9079 N$18158 N$18157 "Straight Waveguide" sch_x=-253 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9080 N$18160 N$18159 "Straight Waveguide" sch_x=-253 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9081 N$18162 N$18161 "Straight Waveguide" sch_x=-253 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9082 N$18164 N$18163 "Straight Waveguide" sch_x=-253 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9083 N$18166 N$18165 "Straight Waveguide" sch_x=-253 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9084 N$18168 N$18167 "Straight Waveguide" sch_x=-253 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9085 N$18170 N$18169 "Straight Waveguide" sch_x=-253 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9086 N$18172 N$18171 "Straight Waveguide" sch_x=-253 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9087 N$18174 N$18173 "Straight Waveguide" sch_x=-251 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9088 N$18176 N$18175 "Straight Waveguide" sch_x=-251 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9089 N$18178 N$18177 "Straight Waveguide" sch_x=-251 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9090 N$18180 N$18179 "Straight Waveguide" sch_x=-251 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9091 N$18182 N$18181 "Straight Waveguide" sch_x=-251 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9092 N$18184 N$18183 "Straight Waveguide" sch_x=-251 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9093 N$18186 N$18185 "Straight Waveguide" sch_x=-251 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9094 N$18188 N$18187 "Straight Waveguide" sch_x=-251 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9095 N$18190 N$18189 "Straight Waveguide" sch_x=-251 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9096 N$18192 N$18191 "Straight Waveguide" sch_x=-251 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9097 N$18194 N$18193 "Straight Waveguide" sch_x=-251 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9098 N$18196 N$18195 "Straight Waveguide" sch_x=-251 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9099 N$18198 N$18197 "Straight Waveguide" sch_x=-251 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9100 N$18200 N$18199 "Straight Waveguide" sch_x=-251 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9101 N$18202 N$18201 "Straight Waveguide" sch_x=-251 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9102 N$18204 N$18203 "Straight Waveguide" sch_x=-251 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9103 N$18206 N$18205 "Straight Waveguide" sch_x=-251 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9104 N$18208 N$18207 "Straight Waveguide" sch_x=-251 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9105 N$18210 N$18209 "Straight Waveguide" sch_x=-251 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9106 N$18212 N$18211 "Straight Waveguide" sch_x=-251 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9107 N$18214 N$18213 "Straight Waveguide" sch_x=-251 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9108 N$18216 N$18215 "Straight Waveguide" sch_x=-251 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9109 N$18218 N$18217 "Straight Waveguide" sch_x=-251 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9110 N$18220 N$18219 "Straight Waveguide" sch_x=-251 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9111 N$18222 N$18221 "Straight Waveguide" sch_x=-251 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9112 N$18224 N$18223 "Straight Waveguide" sch_x=-251 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9113 N$18226 N$18225 "Straight Waveguide" sch_x=-251 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9114 N$18228 N$18227 "Straight Waveguide" sch_x=-251 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9115 N$18230 N$18229 "Straight Waveguide" sch_x=-251 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9116 N$18232 N$18231 "Straight Waveguide" sch_x=-251 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9117 N$18234 N$18233 "Straight Waveguide" sch_x=-251 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9118 N$18236 N$18235 "Straight Waveguide" sch_x=-251 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9119 N$18238 N$18237 "Straight Waveguide" sch_x=-251 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9120 N$18240 N$18239 "Straight Waveguide" sch_x=-251 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9121 N$18242 N$18241 "Straight Waveguide" sch_x=-251 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9122 N$18244 N$18243 "Straight Waveguide" sch_x=-251 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9123 N$18246 N$18245 "Straight Waveguide" sch_x=-251 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9124 N$18248 N$18247 "Straight Waveguide" sch_x=-251 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9125 N$18250 N$18249 "Straight Waveguide" sch_x=-251 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9126 N$18252 N$18251 "Straight Waveguide" sch_x=-251 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9127 N$18254 N$18253 "Straight Waveguide" sch_x=-251 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9128 N$18256 N$18255 "Straight Waveguide" sch_x=-251 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9129 N$18258 N$18257 "Straight Waveguide" sch_x=-251 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9130 N$18260 N$18259 "Straight Waveguide" sch_x=-251 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9131 N$18262 N$18261 "Straight Waveguide" sch_x=-251 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9132 N$18264 N$18263 "Straight Waveguide" sch_x=-251 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9133 N$18266 N$18265 "Straight Waveguide" sch_x=-251 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9134 N$18268 N$18267 "Straight Waveguide" sch_x=-251 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9135 N$18270 N$18269 "Straight Waveguide" sch_x=-251 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9136 N$18272 N$18271 "Straight Waveguide" sch_x=-251 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9137 N$18274 N$18273 "Straight Waveguide" sch_x=-251 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9138 N$18276 N$18275 "Straight Waveguide" sch_x=-251 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9139 N$18278 N$18277 "Straight Waveguide" sch_x=-251 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9140 N$18280 N$18279 "Straight Waveguide" sch_x=-251 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9141 N$18282 N$18281 "Straight Waveguide" sch_x=-251 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9142 N$18284 N$18283 "Straight Waveguide" sch_x=-251 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9143 N$18286 N$18285 "Straight Waveguide" sch_x=-251 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9144 N$18288 N$18287 "Straight Waveguide" sch_x=-251 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9145 N$18290 N$18289 "Straight Waveguide" sch_x=-251 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9146 N$18292 N$18291 "Straight Waveguide" sch_x=-251 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9147 N$18294 N$18293 "Straight Waveguide" sch_x=-251 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9148 N$18296 N$18295 "Straight Waveguide" sch_x=-251 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9149 N$18298 N$18297 "Straight Waveguide" sch_x=-251 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9150 N$18300 N$18299 "Straight Waveguide" sch_x=-251 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9151 N$18302 N$18301 "Straight Waveguide" sch_x=-251 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9152 N$18304 N$18303 "Straight Waveguide" sch_x=-251 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9153 N$18306 N$18305 "Straight Waveguide" sch_x=-251 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9154 N$18308 N$18307 "Straight Waveguide" sch_x=-251 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9155 N$18310 N$18309 "Straight Waveguide" sch_x=-251 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9156 N$18312 N$18311 "Straight Waveguide" sch_x=-251 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9157 N$18314 N$18313 "Straight Waveguide" sch_x=-251 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9158 N$18316 N$18315 "Straight Waveguide" sch_x=-251 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9159 N$18318 N$18317 "Straight Waveguide" sch_x=-251 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9160 N$18320 N$18319 "Straight Waveguide" sch_x=-251 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9161 N$18322 N$18321 "Straight Waveguide" sch_x=-251 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9162 N$18324 N$18323 "Straight Waveguide" sch_x=-251 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9163 N$18326 N$18325 "Straight Waveguide" sch_x=-251 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9164 N$18328 N$18327 "Straight Waveguide" sch_x=-251 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9165 N$18330 N$18329 "Straight Waveguide" sch_x=-251 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9166 N$18332 N$18331 "Straight Waveguide" sch_x=-251 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9167 N$18334 N$18333 "Straight Waveguide" sch_x=-251 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9168 N$18336 N$18335 "Straight Waveguide" sch_x=-251 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9169 N$18338 N$18337 "Straight Waveguide" sch_x=-251 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9170 N$18340 N$18339 "Straight Waveguide" sch_x=-251 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9171 N$18342 N$18341 "Straight Waveguide" sch_x=-251 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9172 N$18344 N$18343 "Straight Waveguide" sch_x=-251 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9173 N$18346 N$18345 "Straight Waveguide" sch_x=-251 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9174 N$18348 N$18347 "Straight Waveguide" sch_x=-251 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9175 N$18350 N$18349 "Straight Waveguide" sch_x=-251 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9176 N$18352 N$18351 "Straight Waveguide" sch_x=-251 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9177 N$18354 N$18353 "Straight Waveguide" sch_x=-251 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9178 N$18356 N$18355 "Straight Waveguide" sch_x=-251 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9179 N$18358 N$18357 "Straight Waveguide" sch_x=-251 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9180 N$18360 N$18359 "Straight Waveguide" sch_x=-251 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9181 N$18362 N$18361 "Straight Waveguide" sch_x=-251 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9182 N$18364 N$18363 "Straight Waveguide" sch_x=-251 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9183 N$18366 N$18365 "Straight Waveguide" sch_x=-251 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9184 N$18368 N$18367 "Straight Waveguide" sch_x=-251 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9185 N$18370 N$18369 "Straight Waveguide" sch_x=-251 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9186 N$18372 N$18371 "Straight Waveguide" sch_x=-251 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9187 N$18374 N$18373 "Straight Waveguide" sch_x=-251 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9188 N$18376 N$18375 "Straight Waveguide" sch_x=-251 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9189 N$18378 N$18377 "Straight Waveguide" sch_x=-251 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9190 N$18380 N$18379 "Straight Waveguide" sch_x=-251 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9191 N$18382 N$18381 "Straight Waveguide" sch_x=-251 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9192 N$18384 N$18383 "Straight Waveguide" sch_x=-251 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9193 N$18386 N$18385 "Straight Waveguide" sch_x=-251 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9194 N$18388 N$18387 "Straight Waveguide" sch_x=-251 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9195 N$18390 N$18389 "Straight Waveguide" sch_x=-251 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9196 N$18392 N$18391 "Straight Waveguide" sch_x=-251 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9197 N$18394 N$18393 "Straight Waveguide" sch_x=-251 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9198 N$18396 N$18395 "Straight Waveguide" sch_x=-251 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9199 N$18398 N$18397 "Straight Waveguide" sch_x=-251 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9200 N$18400 N$18399 "Straight Waveguide" sch_x=-251 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9201 N$18402 N$18401 "Straight Waveguide" sch_x=-251 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9202 N$18404 N$18403 "Straight Waveguide" sch_x=-251 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9203 N$18406 N$18405 "Straight Waveguide" sch_x=-251 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9204 N$18408 N$18407 "Straight Waveguide" sch_x=-251 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9205 N$18410 N$18409 "Straight Waveguide" sch_x=-251 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9206 N$18412 N$18411 "Straight Waveguide" sch_x=-251 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9207 N$18414 N$18413 "Straight Waveguide" sch_x=-251 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9208 N$18416 N$18415 "Straight Waveguide" sch_x=-251 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9209 N$18418 N$18417 "Straight Waveguide" sch_x=-251 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9210 N$18420 N$18419 "Straight Waveguide" sch_x=-251 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9211 N$18422 N$18421 "Straight Waveguide" sch_x=-249 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9212 N$18424 N$18423 "Straight Waveguide" sch_x=-249 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9213 N$18426 N$18425 "Straight Waveguide" sch_x=-249 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9214 N$18428 N$18427 "Straight Waveguide" sch_x=-249 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9215 N$18430 N$18429 "Straight Waveguide" sch_x=-249 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9216 N$18432 N$18431 "Straight Waveguide" sch_x=-249 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9217 N$18434 N$18433 "Straight Waveguide" sch_x=-249 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9218 N$18436 N$18435 "Straight Waveguide" sch_x=-249 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9219 N$18438 N$18437 "Straight Waveguide" sch_x=-249 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9220 N$18440 N$18439 "Straight Waveguide" sch_x=-249 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9221 N$18442 N$18441 "Straight Waveguide" sch_x=-249 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9222 N$18444 N$18443 "Straight Waveguide" sch_x=-249 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9223 N$18446 N$18445 "Straight Waveguide" sch_x=-249 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9224 N$18448 N$18447 "Straight Waveguide" sch_x=-249 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9225 N$18450 N$18449 "Straight Waveguide" sch_x=-249 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9226 N$18452 N$18451 "Straight Waveguide" sch_x=-249 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9227 N$18454 N$18453 "Straight Waveguide" sch_x=-249 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9228 N$18456 N$18455 "Straight Waveguide" sch_x=-249 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9229 N$18458 N$18457 "Straight Waveguide" sch_x=-249 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9230 N$18460 N$18459 "Straight Waveguide" sch_x=-249 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9231 N$18462 N$18461 "Straight Waveguide" sch_x=-249 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9232 N$18464 N$18463 "Straight Waveguide" sch_x=-249 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9233 N$18466 N$18465 "Straight Waveguide" sch_x=-249 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9234 N$18468 N$18467 "Straight Waveguide" sch_x=-249 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9235 N$18470 N$18469 "Straight Waveguide" sch_x=-249 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9236 N$18472 N$18471 "Straight Waveguide" sch_x=-249 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9237 N$18474 N$18473 "Straight Waveguide" sch_x=-249 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9238 N$18476 N$18475 "Straight Waveguide" sch_x=-249 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9239 N$18478 N$18477 "Straight Waveguide" sch_x=-249 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9240 N$18480 N$18479 "Straight Waveguide" sch_x=-249 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9241 N$18482 N$18481 "Straight Waveguide" sch_x=-249 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9242 N$18484 N$18483 "Straight Waveguide" sch_x=-249 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9243 N$18486 N$18485 "Straight Waveguide" sch_x=-249 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9244 N$18488 N$18487 "Straight Waveguide" sch_x=-249 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9245 N$18490 N$18489 "Straight Waveguide" sch_x=-249 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9246 N$18492 N$18491 "Straight Waveguide" sch_x=-249 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9247 N$18494 N$18493 "Straight Waveguide" sch_x=-249 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9248 N$18496 N$18495 "Straight Waveguide" sch_x=-249 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9249 N$18498 N$18497 "Straight Waveguide" sch_x=-249 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9250 N$18500 N$18499 "Straight Waveguide" sch_x=-249 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9251 N$18502 N$18501 "Straight Waveguide" sch_x=-249 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9252 N$18504 N$18503 "Straight Waveguide" sch_x=-249 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9253 N$18506 N$18505 "Straight Waveguide" sch_x=-249 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9254 N$18508 N$18507 "Straight Waveguide" sch_x=-249 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9255 N$18510 N$18509 "Straight Waveguide" sch_x=-249 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9256 N$18512 N$18511 "Straight Waveguide" sch_x=-249 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9257 N$18514 N$18513 "Straight Waveguide" sch_x=-249 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9258 N$18516 N$18515 "Straight Waveguide" sch_x=-249 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9259 N$18518 N$18517 "Straight Waveguide" sch_x=-249 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9260 N$18520 N$18519 "Straight Waveguide" sch_x=-249 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9261 N$18522 N$18521 "Straight Waveguide" sch_x=-249 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9262 N$18524 N$18523 "Straight Waveguide" sch_x=-249 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9263 N$18526 N$18525 "Straight Waveguide" sch_x=-249 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9264 N$18528 N$18527 "Straight Waveguide" sch_x=-249 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9265 N$18530 N$18529 "Straight Waveguide" sch_x=-249 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9266 N$18532 N$18531 "Straight Waveguide" sch_x=-249 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9267 N$18534 N$18533 "Straight Waveguide" sch_x=-249 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9268 N$18536 N$18535 "Straight Waveguide" sch_x=-249 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9269 N$18538 N$18537 "Straight Waveguide" sch_x=-249 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9270 N$18540 N$18539 "Straight Waveguide" sch_x=-249 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9271 N$18542 N$18541 "Straight Waveguide" sch_x=-249 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9272 N$18544 N$18543 "Straight Waveguide" sch_x=-249 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9273 N$18546 N$18545 "Straight Waveguide" sch_x=-249 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9274 N$18548 N$18547 "Straight Waveguide" sch_x=-249 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9275 N$18550 N$18549 "Straight Waveguide" sch_x=-249 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9276 N$18552 N$18551 "Straight Waveguide" sch_x=-249 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9277 N$18554 N$18553 "Straight Waveguide" sch_x=-249 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9278 N$18556 N$18555 "Straight Waveguide" sch_x=-249 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9279 N$18558 N$18557 "Straight Waveguide" sch_x=-249 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9280 N$18560 N$18559 "Straight Waveguide" sch_x=-249 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9281 N$18562 N$18561 "Straight Waveguide" sch_x=-249 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9282 N$18564 N$18563 "Straight Waveguide" sch_x=-249 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9283 N$18566 N$18565 "Straight Waveguide" sch_x=-249 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9284 N$18568 N$18567 "Straight Waveguide" sch_x=-249 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9285 N$18570 N$18569 "Straight Waveguide" sch_x=-249 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9286 N$18572 N$18571 "Straight Waveguide" sch_x=-249 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9287 N$18574 N$18573 "Straight Waveguide" sch_x=-249 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9288 N$18576 N$18575 "Straight Waveguide" sch_x=-249 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9289 N$18578 N$18577 "Straight Waveguide" sch_x=-249 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9290 N$18580 N$18579 "Straight Waveguide" sch_x=-249 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9291 N$18582 N$18581 "Straight Waveguide" sch_x=-249 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9292 N$18584 N$18583 "Straight Waveguide" sch_x=-249 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9293 N$18586 N$18585 "Straight Waveguide" sch_x=-249 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9294 N$18588 N$18587 "Straight Waveguide" sch_x=-249 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9295 N$18590 N$18589 "Straight Waveguide" sch_x=-249 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9296 N$18592 N$18591 "Straight Waveguide" sch_x=-249 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9297 N$18594 N$18593 "Straight Waveguide" sch_x=-249 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9298 N$18596 N$18595 "Straight Waveguide" sch_x=-249 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9299 N$18598 N$18597 "Straight Waveguide" sch_x=-249 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9300 N$18600 N$18599 "Straight Waveguide" sch_x=-249 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9301 N$18602 N$18601 "Straight Waveguide" sch_x=-249 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9302 N$18604 N$18603 "Straight Waveguide" sch_x=-249 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9303 N$18606 N$18605 "Straight Waveguide" sch_x=-249 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9304 N$18608 N$18607 "Straight Waveguide" sch_x=-249 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9305 N$18610 N$18609 "Straight Waveguide" sch_x=-249 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9306 N$18612 N$18611 "Straight Waveguide" sch_x=-249 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9307 N$18614 N$18613 "Straight Waveguide" sch_x=-249 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9308 N$18616 N$18615 "Straight Waveguide" sch_x=-249 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9309 N$18618 N$18617 "Straight Waveguide" sch_x=-249 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9310 N$18620 N$18619 "Straight Waveguide" sch_x=-249 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9311 N$18622 N$18621 "Straight Waveguide" sch_x=-249 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9312 N$18624 N$18623 "Straight Waveguide" sch_x=-249 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9313 N$18626 N$18625 "Straight Waveguide" sch_x=-249 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9314 N$18628 N$18627 "Straight Waveguide" sch_x=-249 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9315 N$18630 N$18629 "Straight Waveguide" sch_x=-249 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9316 N$18632 N$18631 "Straight Waveguide" sch_x=-249 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9317 N$18634 N$18633 "Straight Waveguide" sch_x=-249 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9318 N$18636 N$18635 "Straight Waveguide" sch_x=-249 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9319 N$18638 N$18637 "Straight Waveguide" sch_x=-249 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9320 N$18640 N$18639 "Straight Waveguide" sch_x=-249 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9321 N$18642 N$18641 "Straight Waveguide" sch_x=-249 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9322 N$18644 N$18643 "Straight Waveguide" sch_x=-249 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9323 N$18646 N$18645 "Straight Waveguide" sch_x=-249 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9324 N$18648 N$18647 "Straight Waveguide" sch_x=-249 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9325 N$18650 N$18649 "Straight Waveguide" sch_x=-249 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9326 N$18652 N$18651 "Straight Waveguide" sch_x=-249 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9327 N$18654 N$18653 "Straight Waveguide" sch_x=-249 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9328 N$18656 N$18655 "Straight Waveguide" sch_x=-249 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9329 N$18658 N$18657 "Straight Waveguide" sch_x=-249 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9330 N$18660 N$18659 "Straight Waveguide" sch_x=-249 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9331 N$18662 N$18661 "Straight Waveguide" sch_x=-249 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9332 N$18664 N$18663 "Straight Waveguide" sch_x=-249 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9333 N$18666 N$18665 "Straight Waveguide" sch_x=-247 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9334 N$18668 N$18667 "Straight Waveguide" sch_x=-247 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9335 N$18670 N$18669 "Straight Waveguide" sch_x=-247 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9336 N$18672 N$18671 "Straight Waveguide" sch_x=-247 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9337 N$18674 N$18673 "Straight Waveguide" sch_x=-247 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9338 N$18676 N$18675 "Straight Waveguide" sch_x=-247 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9339 N$18678 N$18677 "Straight Waveguide" sch_x=-247 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9340 N$18680 N$18679 "Straight Waveguide" sch_x=-247 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9341 N$18682 N$18681 "Straight Waveguide" sch_x=-247 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9342 N$18684 N$18683 "Straight Waveguide" sch_x=-247 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9343 N$18686 N$18685 "Straight Waveguide" sch_x=-247 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9344 N$18688 N$18687 "Straight Waveguide" sch_x=-247 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9345 N$18690 N$18689 "Straight Waveguide" sch_x=-247 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9346 N$18692 N$18691 "Straight Waveguide" sch_x=-247 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9347 N$18694 N$18693 "Straight Waveguide" sch_x=-247 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9348 N$18696 N$18695 "Straight Waveguide" sch_x=-247 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9349 N$18698 N$18697 "Straight Waveguide" sch_x=-247 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9350 N$18700 N$18699 "Straight Waveguide" sch_x=-247 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9351 N$18702 N$18701 "Straight Waveguide" sch_x=-247 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9352 N$18704 N$18703 "Straight Waveguide" sch_x=-247 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9353 N$18706 N$18705 "Straight Waveguide" sch_x=-247 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9354 N$18708 N$18707 "Straight Waveguide" sch_x=-247 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9355 N$18710 N$18709 "Straight Waveguide" sch_x=-247 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9356 N$18712 N$18711 "Straight Waveguide" sch_x=-247 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9357 N$18714 N$18713 "Straight Waveguide" sch_x=-247 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9358 N$18716 N$18715 "Straight Waveguide" sch_x=-247 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9359 N$18718 N$18717 "Straight Waveguide" sch_x=-247 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9360 N$18720 N$18719 "Straight Waveguide" sch_x=-247 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9361 N$18722 N$18721 "Straight Waveguide" sch_x=-247 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9362 N$18724 N$18723 "Straight Waveguide" sch_x=-247 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9363 N$18726 N$18725 "Straight Waveguide" sch_x=-247 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9364 N$18728 N$18727 "Straight Waveguide" sch_x=-247 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9365 N$18730 N$18729 "Straight Waveguide" sch_x=-247 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9366 N$18732 N$18731 "Straight Waveguide" sch_x=-247 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9367 N$18734 N$18733 "Straight Waveguide" sch_x=-247 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9368 N$18736 N$18735 "Straight Waveguide" sch_x=-247 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9369 N$18738 N$18737 "Straight Waveguide" sch_x=-247 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9370 N$18740 N$18739 "Straight Waveguide" sch_x=-247 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9371 N$18742 N$18741 "Straight Waveguide" sch_x=-247 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9372 N$18744 N$18743 "Straight Waveguide" sch_x=-247 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9373 N$18746 N$18745 "Straight Waveguide" sch_x=-247 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9374 N$18748 N$18747 "Straight Waveguide" sch_x=-247 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9375 N$18750 N$18749 "Straight Waveguide" sch_x=-247 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9376 N$18752 N$18751 "Straight Waveguide" sch_x=-247 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9377 N$18754 N$18753 "Straight Waveguide" sch_x=-247 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9378 N$18756 N$18755 "Straight Waveguide" sch_x=-247 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9379 N$18758 N$18757 "Straight Waveguide" sch_x=-247 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9380 N$18760 N$18759 "Straight Waveguide" sch_x=-247 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9381 N$18762 N$18761 "Straight Waveguide" sch_x=-247 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9382 N$18764 N$18763 "Straight Waveguide" sch_x=-247 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9383 N$18766 N$18765 "Straight Waveguide" sch_x=-247 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9384 N$18768 N$18767 "Straight Waveguide" sch_x=-247 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9385 N$18770 N$18769 "Straight Waveguide" sch_x=-247 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9386 N$18772 N$18771 "Straight Waveguide" sch_x=-247 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9387 N$18774 N$18773 "Straight Waveguide" sch_x=-247 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9388 N$18776 N$18775 "Straight Waveguide" sch_x=-247 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9389 N$18778 N$18777 "Straight Waveguide" sch_x=-247 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9390 N$18780 N$18779 "Straight Waveguide" sch_x=-247 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9391 N$18782 N$18781 "Straight Waveguide" sch_x=-247 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9392 N$18784 N$18783 "Straight Waveguide" sch_x=-247 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9393 N$18786 N$18785 "Straight Waveguide" sch_x=-247 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9394 N$18788 N$18787 "Straight Waveguide" sch_x=-247 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9395 N$18790 N$18789 "Straight Waveguide" sch_x=-247 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9396 N$18792 N$18791 "Straight Waveguide" sch_x=-247 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9397 N$18794 N$18793 "Straight Waveguide" sch_x=-247 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9398 N$18796 N$18795 "Straight Waveguide" sch_x=-247 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9399 N$18798 N$18797 "Straight Waveguide" sch_x=-247 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9400 N$18800 N$18799 "Straight Waveguide" sch_x=-247 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9401 N$18802 N$18801 "Straight Waveguide" sch_x=-247 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9402 N$18804 N$18803 "Straight Waveguide" sch_x=-247 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9403 N$18806 N$18805 "Straight Waveguide" sch_x=-247 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9404 N$18808 N$18807 "Straight Waveguide" sch_x=-247 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9405 N$18810 N$18809 "Straight Waveguide" sch_x=-247 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9406 N$18812 N$18811 "Straight Waveguide" sch_x=-247 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9407 N$18814 N$18813 "Straight Waveguide" sch_x=-247 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9408 N$18816 N$18815 "Straight Waveguide" sch_x=-247 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9409 N$18818 N$18817 "Straight Waveguide" sch_x=-247 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9410 N$18820 N$18819 "Straight Waveguide" sch_x=-247 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9411 N$18822 N$18821 "Straight Waveguide" sch_x=-247 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9412 N$18824 N$18823 "Straight Waveguide" sch_x=-247 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9413 N$18826 N$18825 "Straight Waveguide" sch_x=-247 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9414 N$18828 N$18827 "Straight Waveguide" sch_x=-247 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9415 N$18830 N$18829 "Straight Waveguide" sch_x=-247 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9416 N$18832 N$18831 "Straight Waveguide" sch_x=-247 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9417 N$18834 N$18833 "Straight Waveguide" sch_x=-247 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9418 N$18836 N$18835 "Straight Waveguide" sch_x=-247 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9419 N$18838 N$18837 "Straight Waveguide" sch_x=-247 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9420 N$18840 N$18839 "Straight Waveguide" sch_x=-247 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9421 N$18842 N$18841 "Straight Waveguide" sch_x=-247 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9422 N$18844 N$18843 "Straight Waveguide" sch_x=-247 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9423 N$18846 N$18845 "Straight Waveguide" sch_x=-247 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9424 N$18848 N$18847 "Straight Waveguide" sch_x=-247 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9425 N$18850 N$18849 "Straight Waveguide" sch_x=-247 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9426 N$18852 N$18851 "Straight Waveguide" sch_x=-247 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9427 N$18854 N$18853 "Straight Waveguide" sch_x=-247 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9428 N$18856 N$18855 "Straight Waveguide" sch_x=-247 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9429 N$18858 N$18857 "Straight Waveguide" sch_x=-247 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9430 N$18860 N$18859 "Straight Waveguide" sch_x=-247 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9431 N$18862 N$18861 "Straight Waveguide" sch_x=-247 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9432 N$18864 N$18863 "Straight Waveguide" sch_x=-247 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9433 N$18866 N$18865 "Straight Waveguide" sch_x=-247 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9434 N$18868 N$18867 "Straight Waveguide" sch_x=-247 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9435 N$18870 N$18869 "Straight Waveguide" sch_x=-247 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9436 N$18872 N$18871 "Straight Waveguide" sch_x=-247 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9437 N$18874 N$18873 "Straight Waveguide" sch_x=-247 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9438 N$18876 N$18875 "Straight Waveguide" sch_x=-247 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9439 N$18878 N$18877 "Straight Waveguide" sch_x=-247 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9440 N$18880 N$18879 "Straight Waveguide" sch_x=-247 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9441 N$18882 N$18881 "Straight Waveguide" sch_x=-247 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9442 N$18884 N$18883 "Straight Waveguide" sch_x=-247 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9443 N$18886 N$18885 "Straight Waveguide" sch_x=-247 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9444 N$18888 N$18887 "Straight Waveguide" sch_x=-247 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9445 N$18890 N$18889 "Straight Waveguide" sch_x=-247 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9446 N$18892 N$18891 "Straight Waveguide" sch_x=-247 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9447 N$18894 N$18893 "Straight Waveguide" sch_x=-247 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9448 N$18896 N$18895 "Straight Waveguide" sch_x=-247 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9449 N$18898 N$18897 "Straight Waveguide" sch_x=-247 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9450 N$18900 N$18899 "Straight Waveguide" sch_x=-247 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9451 N$18902 N$18901 "Straight Waveguide" sch_x=-247 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9452 N$18904 N$18903 "Straight Waveguide" sch_x=-247 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9453 N$18906 N$18905 "Straight Waveguide" sch_x=-245 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9454 N$18908 N$18907 "Straight Waveguide" sch_x=-245 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9455 N$18910 N$18909 "Straight Waveguide" sch_x=-245 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9456 N$18912 N$18911 "Straight Waveguide" sch_x=-245 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9457 N$18914 N$18913 "Straight Waveguide" sch_x=-245 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9458 N$18916 N$18915 "Straight Waveguide" sch_x=-245 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9459 N$18918 N$18917 "Straight Waveguide" sch_x=-245 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9460 N$18920 N$18919 "Straight Waveguide" sch_x=-245 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9461 N$18922 N$18921 "Straight Waveguide" sch_x=-245 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9462 N$18924 N$18923 "Straight Waveguide" sch_x=-245 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9463 N$18926 N$18925 "Straight Waveguide" sch_x=-245 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9464 N$18928 N$18927 "Straight Waveguide" sch_x=-245 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9465 N$18930 N$18929 "Straight Waveguide" sch_x=-245 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9466 N$18932 N$18931 "Straight Waveguide" sch_x=-245 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9467 N$18934 N$18933 "Straight Waveguide" sch_x=-245 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9468 N$18936 N$18935 "Straight Waveguide" sch_x=-245 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9469 N$18938 N$18937 "Straight Waveguide" sch_x=-245 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9470 N$18940 N$18939 "Straight Waveguide" sch_x=-245 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9471 N$18942 N$18941 "Straight Waveguide" sch_x=-245 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9472 N$18944 N$18943 "Straight Waveguide" sch_x=-245 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9473 N$18946 N$18945 "Straight Waveguide" sch_x=-245 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9474 N$18948 N$18947 "Straight Waveguide" sch_x=-245 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9475 N$18950 N$18949 "Straight Waveguide" sch_x=-245 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9476 N$18952 N$18951 "Straight Waveguide" sch_x=-245 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9477 N$18954 N$18953 "Straight Waveguide" sch_x=-245 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9478 N$18956 N$18955 "Straight Waveguide" sch_x=-245 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9479 N$18958 N$18957 "Straight Waveguide" sch_x=-245 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9480 N$18960 N$18959 "Straight Waveguide" sch_x=-245 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9481 N$18962 N$18961 "Straight Waveguide" sch_x=-245 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9482 N$18964 N$18963 "Straight Waveguide" sch_x=-245 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9483 N$18966 N$18965 "Straight Waveguide" sch_x=-245 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9484 N$18968 N$18967 "Straight Waveguide" sch_x=-245 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9485 N$18970 N$18969 "Straight Waveguide" sch_x=-245 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9486 N$18972 N$18971 "Straight Waveguide" sch_x=-245 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9487 N$18974 N$18973 "Straight Waveguide" sch_x=-245 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9488 N$18976 N$18975 "Straight Waveguide" sch_x=-245 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9489 N$18978 N$18977 "Straight Waveguide" sch_x=-245 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9490 N$18980 N$18979 "Straight Waveguide" sch_x=-245 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9491 N$18982 N$18981 "Straight Waveguide" sch_x=-245 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9492 N$18984 N$18983 "Straight Waveguide" sch_x=-245 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9493 N$18986 N$18985 "Straight Waveguide" sch_x=-245 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9494 N$18988 N$18987 "Straight Waveguide" sch_x=-245 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9495 N$18990 N$18989 "Straight Waveguide" sch_x=-245 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9496 N$18992 N$18991 "Straight Waveguide" sch_x=-245 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9497 N$18994 N$18993 "Straight Waveguide" sch_x=-245 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9498 N$18996 N$18995 "Straight Waveguide" sch_x=-245 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9499 N$18998 N$18997 "Straight Waveguide" sch_x=-245 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9500 N$19000 N$18999 "Straight Waveguide" sch_x=-245 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9501 N$19002 N$19001 "Straight Waveguide" sch_x=-245 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9502 N$19004 N$19003 "Straight Waveguide" sch_x=-245 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9503 N$19006 N$19005 "Straight Waveguide" sch_x=-245 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9504 N$19008 N$19007 "Straight Waveguide" sch_x=-245 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9505 N$19010 N$19009 "Straight Waveguide" sch_x=-245 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9506 N$19012 N$19011 "Straight Waveguide" sch_x=-245 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9507 N$19014 N$19013 "Straight Waveguide" sch_x=-245 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9508 N$19016 N$19015 "Straight Waveguide" sch_x=-245 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9509 N$19018 N$19017 "Straight Waveguide" sch_x=-245 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9510 N$19020 N$19019 "Straight Waveguide" sch_x=-245 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9511 N$19022 N$19021 "Straight Waveguide" sch_x=-245 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9512 N$19024 N$19023 "Straight Waveguide" sch_x=-245 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9513 N$19026 N$19025 "Straight Waveguide" sch_x=-245 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9514 N$19028 N$19027 "Straight Waveguide" sch_x=-245 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9515 N$19030 N$19029 "Straight Waveguide" sch_x=-245 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9516 N$19032 N$19031 "Straight Waveguide" sch_x=-245 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9517 N$19034 N$19033 "Straight Waveguide" sch_x=-245 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9518 N$19036 N$19035 "Straight Waveguide" sch_x=-245 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9519 N$19038 N$19037 "Straight Waveguide" sch_x=-245 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9520 N$19040 N$19039 "Straight Waveguide" sch_x=-245 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9521 N$19042 N$19041 "Straight Waveguide" sch_x=-245 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9522 N$19044 N$19043 "Straight Waveguide" sch_x=-245 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9523 N$19046 N$19045 "Straight Waveguide" sch_x=-245 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9524 N$19048 N$19047 "Straight Waveguide" sch_x=-245 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9525 N$19050 N$19049 "Straight Waveguide" sch_x=-245 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9526 N$19052 N$19051 "Straight Waveguide" sch_x=-245 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9527 N$19054 N$19053 "Straight Waveguide" sch_x=-245 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9528 N$19056 N$19055 "Straight Waveguide" sch_x=-245 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9529 N$19058 N$19057 "Straight Waveguide" sch_x=-245 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9530 N$19060 N$19059 "Straight Waveguide" sch_x=-245 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9531 N$19062 N$19061 "Straight Waveguide" sch_x=-245 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9532 N$19064 N$19063 "Straight Waveguide" sch_x=-245 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9533 N$19066 N$19065 "Straight Waveguide" sch_x=-245 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9534 N$19068 N$19067 "Straight Waveguide" sch_x=-245 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9535 N$19070 N$19069 "Straight Waveguide" sch_x=-245 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9536 N$19072 N$19071 "Straight Waveguide" sch_x=-245 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9537 N$19074 N$19073 "Straight Waveguide" sch_x=-245 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9538 N$19076 N$19075 "Straight Waveguide" sch_x=-245 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9539 N$19078 N$19077 "Straight Waveguide" sch_x=-245 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9540 N$19080 N$19079 "Straight Waveguide" sch_x=-245 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9541 N$19082 N$19081 "Straight Waveguide" sch_x=-245 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9542 N$19084 N$19083 "Straight Waveguide" sch_x=-245 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9543 N$19086 N$19085 "Straight Waveguide" sch_x=-245 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9544 N$19088 N$19087 "Straight Waveguide" sch_x=-245 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9545 N$19090 N$19089 "Straight Waveguide" sch_x=-245 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9546 N$19092 N$19091 "Straight Waveguide" sch_x=-245 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9547 N$19094 N$19093 "Straight Waveguide" sch_x=-245 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9548 N$19096 N$19095 "Straight Waveguide" sch_x=-245 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9549 N$19098 N$19097 "Straight Waveguide" sch_x=-245 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9550 N$19100 N$19099 "Straight Waveguide" sch_x=-245 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9551 N$19102 N$19101 "Straight Waveguide" sch_x=-245 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9552 N$19104 N$19103 "Straight Waveguide" sch_x=-245 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9553 N$19106 N$19105 "Straight Waveguide" sch_x=-245 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9554 N$19108 N$19107 "Straight Waveguide" sch_x=-245 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9555 N$19110 N$19109 "Straight Waveguide" sch_x=-245 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9556 N$19112 N$19111 "Straight Waveguide" sch_x=-245 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9557 N$19114 N$19113 "Straight Waveguide" sch_x=-245 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9558 N$19116 N$19115 "Straight Waveguide" sch_x=-245 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9559 N$19118 N$19117 "Straight Waveguide" sch_x=-245 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9560 N$19120 N$19119 "Straight Waveguide" sch_x=-245 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9561 N$19122 N$19121 "Straight Waveguide" sch_x=-245 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9562 N$19124 N$19123 "Straight Waveguide" sch_x=-245 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9563 N$19126 N$19125 "Straight Waveguide" sch_x=-245 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9564 N$19128 N$19127 "Straight Waveguide" sch_x=-245 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9565 N$19130 N$19129 "Straight Waveguide" sch_x=-245 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9566 N$19132 N$19131 "Straight Waveguide" sch_x=-245 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9567 N$19134 N$19133 "Straight Waveguide" sch_x=-245 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9568 N$19136 N$19135 "Straight Waveguide" sch_x=-245 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9569 N$19138 N$19137 "Straight Waveguide" sch_x=-245 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9570 N$19140 N$19139 "Straight Waveguide" sch_x=-245 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9571 N$19142 N$19141 "Straight Waveguide" sch_x=-243 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9572 N$19144 N$19143 "Straight Waveguide" sch_x=-243 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9573 N$19146 N$19145 "Straight Waveguide" sch_x=-243 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9574 N$19148 N$19147 "Straight Waveguide" sch_x=-243 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9575 N$19150 N$19149 "Straight Waveguide" sch_x=-243 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9576 N$19152 N$19151 "Straight Waveguide" sch_x=-243 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9577 N$19154 N$19153 "Straight Waveguide" sch_x=-243 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9578 N$19156 N$19155 "Straight Waveguide" sch_x=-243 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9579 N$19158 N$19157 "Straight Waveguide" sch_x=-243 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9580 N$19160 N$19159 "Straight Waveguide" sch_x=-243 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9581 N$19162 N$19161 "Straight Waveguide" sch_x=-243 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9582 N$19164 N$19163 "Straight Waveguide" sch_x=-243 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9583 N$19166 N$19165 "Straight Waveguide" sch_x=-243 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9584 N$19168 N$19167 "Straight Waveguide" sch_x=-243 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9585 N$19170 N$19169 "Straight Waveguide" sch_x=-243 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9586 N$19172 N$19171 "Straight Waveguide" sch_x=-243 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9587 N$19174 N$19173 "Straight Waveguide" sch_x=-243 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9588 N$19176 N$19175 "Straight Waveguide" sch_x=-243 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9589 N$19178 N$19177 "Straight Waveguide" sch_x=-243 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9590 N$19180 N$19179 "Straight Waveguide" sch_x=-243 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9591 N$19182 N$19181 "Straight Waveguide" sch_x=-243 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9592 N$19184 N$19183 "Straight Waveguide" sch_x=-243 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9593 N$19186 N$19185 "Straight Waveguide" sch_x=-243 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9594 N$19188 N$19187 "Straight Waveguide" sch_x=-243 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9595 N$19190 N$19189 "Straight Waveguide" sch_x=-243 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9596 N$19192 N$19191 "Straight Waveguide" sch_x=-243 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9597 N$19194 N$19193 "Straight Waveguide" sch_x=-243 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9598 N$19196 N$19195 "Straight Waveguide" sch_x=-243 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9599 N$19198 N$19197 "Straight Waveguide" sch_x=-243 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9600 N$19200 N$19199 "Straight Waveguide" sch_x=-243 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9601 N$19202 N$19201 "Straight Waveguide" sch_x=-243 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9602 N$19204 N$19203 "Straight Waveguide" sch_x=-243 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9603 N$19206 N$19205 "Straight Waveguide" sch_x=-243 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9604 N$19208 N$19207 "Straight Waveguide" sch_x=-243 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9605 N$19210 N$19209 "Straight Waveguide" sch_x=-243 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9606 N$19212 N$19211 "Straight Waveguide" sch_x=-243 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9607 N$19214 N$19213 "Straight Waveguide" sch_x=-243 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9608 N$19216 N$19215 "Straight Waveguide" sch_x=-243 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9609 N$19218 N$19217 "Straight Waveguide" sch_x=-243 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9610 N$19220 N$19219 "Straight Waveguide" sch_x=-243 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9611 N$19222 N$19221 "Straight Waveguide" sch_x=-243 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9612 N$19224 N$19223 "Straight Waveguide" sch_x=-243 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9613 N$19226 N$19225 "Straight Waveguide" sch_x=-243 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9614 N$19228 N$19227 "Straight Waveguide" sch_x=-243 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9615 N$19230 N$19229 "Straight Waveguide" sch_x=-243 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9616 N$19232 N$19231 "Straight Waveguide" sch_x=-243 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9617 N$19234 N$19233 "Straight Waveguide" sch_x=-243 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9618 N$19236 N$19235 "Straight Waveguide" sch_x=-243 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9619 N$19238 N$19237 "Straight Waveguide" sch_x=-243 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9620 N$19240 N$19239 "Straight Waveguide" sch_x=-243 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9621 N$19242 N$19241 "Straight Waveguide" sch_x=-243 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9622 N$19244 N$19243 "Straight Waveguide" sch_x=-243 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9623 N$19246 N$19245 "Straight Waveguide" sch_x=-243 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9624 N$19248 N$19247 "Straight Waveguide" sch_x=-243 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9625 N$19250 N$19249 "Straight Waveguide" sch_x=-243 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9626 N$19252 N$19251 "Straight Waveguide" sch_x=-243 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9627 N$19254 N$19253 "Straight Waveguide" sch_x=-243 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9628 N$19256 N$19255 "Straight Waveguide" sch_x=-243 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9629 N$19258 N$19257 "Straight Waveguide" sch_x=-243 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9630 N$19260 N$19259 "Straight Waveguide" sch_x=-243 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9631 N$19262 N$19261 "Straight Waveguide" sch_x=-243 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9632 N$19264 N$19263 "Straight Waveguide" sch_x=-243 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9633 N$19266 N$19265 "Straight Waveguide" sch_x=-243 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9634 N$19268 N$19267 "Straight Waveguide" sch_x=-243 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9635 N$19270 N$19269 "Straight Waveguide" sch_x=-243 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9636 N$19272 N$19271 "Straight Waveguide" sch_x=-243 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9637 N$19274 N$19273 "Straight Waveguide" sch_x=-243 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9638 N$19276 N$19275 "Straight Waveguide" sch_x=-243 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9639 N$19278 N$19277 "Straight Waveguide" sch_x=-243 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9640 N$19280 N$19279 "Straight Waveguide" sch_x=-243 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9641 N$19282 N$19281 "Straight Waveguide" sch_x=-243 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9642 N$19284 N$19283 "Straight Waveguide" sch_x=-243 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9643 N$19286 N$19285 "Straight Waveguide" sch_x=-243 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9644 N$19288 N$19287 "Straight Waveguide" sch_x=-243 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9645 N$19290 N$19289 "Straight Waveguide" sch_x=-243 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9646 N$19292 N$19291 "Straight Waveguide" sch_x=-243 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9647 N$19294 N$19293 "Straight Waveguide" sch_x=-243 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9648 N$19296 N$19295 "Straight Waveguide" sch_x=-243 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9649 N$19298 N$19297 "Straight Waveguide" sch_x=-243 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9650 N$19300 N$19299 "Straight Waveguide" sch_x=-243 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9651 N$19302 N$19301 "Straight Waveguide" sch_x=-243 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9652 N$19304 N$19303 "Straight Waveguide" sch_x=-243 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9653 N$19306 N$19305 "Straight Waveguide" sch_x=-243 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9654 N$19308 N$19307 "Straight Waveguide" sch_x=-243 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9655 N$19310 N$19309 "Straight Waveguide" sch_x=-243 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9656 N$19312 N$19311 "Straight Waveguide" sch_x=-243 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9657 N$19314 N$19313 "Straight Waveguide" sch_x=-243 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9658 N$19316 N$19315 "Straight Waveguide" sch_x=-243 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9659 N$19318 N$19317 "Straight Waveguide" sch_x=-243 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9660 N$19320 N$19319 "Straight Waveguide" sch_x=-243 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9661 N$19322 N$19321 "Straight Waveguide" sch_x=-243 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9662 N$19324 N$19323 "Straight Waveguide" sch_x=-243 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9663 N$19326 N$19325 "Straight Waveguide" sch_x=-243 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9664 N$19328 N$19327 "Straight Waveguide" sch_x=-243 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9665 N$19330 N$19329 "Straight Waveguide" sch_x=-243 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9666 N$19332 N$19331 "Straight Waveguide" sch_x=-243 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9667 N$19334 N$19333 "Straight Waveguide" sch_x=-243 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9668 N$19336 N$19335 "Straight Waveguide" sch_x=-243 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9669 N$19338 N$19337 "Straight Waveguide" sch_x=-243 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9670 N$19340 N$19339 "Straight Waveguide" sch_x=-243 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9671 N$19342 N$19341 "Straight Waveguide" sch_x=-243 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9672 N$19344 N$19343 "Straight Waveguide" sch_x=-243 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9673 N$19346 N$19345 "Straight Waveguide" sch_x=-243 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9674 N$19348 N$19347 "Straight Waveguide" sch_x=-243 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9675 N$19350 N$19349 "Straight Waveguide" sch_x=-243 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9676 N$19352 N$19351 "Straight Waveguide" sch_x=-243 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9677 N$19354 N$19353 "Straight Waveguide" sch_x=-243 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9678 N$19356 N$19355 "Straight Waveguide" sch_x=-243 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9679 N$19358 N$19357 "Straight Waveguide" sch_x=-243 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9680 N$19360 N$19359 "Straight Waveguide" sch_x=-243 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9681 N$19362 N$19361 "Straight Waveguide" sch_x=-243 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9682 N$19364 N$19363 "Straight Waveguide" sch_x=-243 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9683 N$19366 N$19365 "Straight Waveguide" sch_x=-243 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9684 N$19368 N$19367 "Straight Waveguide" sch_x=-243 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9685 N$19370 N$19369 "Straight Waveguide" sch_x=-243 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9686 N$19372 N$19371 "Straight Waveguide" sch_x=-243 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9687 N$19374 N$19373 "Straight Waveguide" sch_x=-241 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9688 N$19376 N$19375 "Straight Waveguide" sch_x=-241 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9689 N$19378 N$19377 "Straight Waveguide" sch_x=-241 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9690 N$19380 N$19379 "Straight Waveguide" sch_x=-241 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9691 N$19382 N$19381 "Straight Waveguide" sch_x=-241 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9692 N$19384 N$19383 "Straight Waveguide" sch_x=-241 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9693 N$19386 N$19385 "Straight Waveguide" sch_x=-241 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9694 N$19388 N$19387 "Straight Waveguide" sch_x=-241 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9695 N$19390 N$19389 "Straight Waveguide" sch_x=-241 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9696 N$19392 N$19391 "Straight Waveguide" sch_x=-241 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9697 N$19394 N$19393 "Straight Waveguide" sch_x=-241 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9698 N$19396 N$19395 "Straight Waveguide" sch_x=-241 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9699 N$19398 N$19397 "Straight Waveguide" sch_x=-241 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9700 N$19400 N$19399 "Straight Waveguide" sch_x=-241 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9701 N$19402 N$19401 "Straight Waveguide" sch_x=-241 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9702 N$19404 N$19403 "Straight Waveguide" sch_x=-241 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9703 N$19406 N$19405 "Straight Waveguide" sch_x=-241 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9704 N$19408 N$19407 "Straight Waveguide" sch_x=-241 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9705 N$19410 N$19409 "Straight Waveguide" sch_x=-241 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9706 N$19412 N$19411 "Straight Waveguide" sch_x=-241 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9707 N$19414 N$19413 "Straight Waveguide" sch_x=-241 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9708 N$19416 N$19415 "Straight Waveguide" sch_x=-241 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9709 N$19418 N$19417 "Straight Waveguide" sch_x=-241 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9710 N$19420 N$19419 "Straight Waveguide" sch_x=-241 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9711 N$19422 N$19421 "Straight Waveguide" sch_x=-241 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9712 N$19424 N$19423 "Straight Waveguide" sch_x=-241 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9713 N$19426 N$19425 "Straight Waveguide" sch_x=-241 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9714 N$19428 N$19427 "Straight Waveguide" sch_x=-241 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9715 N$19430 N$19429 "Straight Waveguide" sch_x=-241 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9716 N$19432 N$19431 "Straight Waveguide" sch_x=-241 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9717 N$19434 N$19433 "Straight Waveguide" sch_x=-241 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9718 N$19436 N$19435 "Straight Waveguide" sch_x=-241 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9719 N$19438 N$19437 "Straight Waveguide" sch_x=-241 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9720 N$19440 N$19439 "Straight Waveguide" sch_x=-241 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9721 N$19442 N$19441 "Straight Waveguide" sch_x=-241 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9722 N$19444 N$19443 "Straight Waveguide" sch_x=-241 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9723 N$19446 N$19445 "Straight Waveguide" sch_x=-241 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9724 N$19448 N$19447 "Straight Waveguide" sch_x=-241 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9725 N$19450 N$19449 "Straight Waveguide" sch_x=-241 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9726 N$19452 N$19451 "Straight Waveguide" sch_x=-241 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9727 N$19454 N$19453 "Straight Waveguide" sch_x=-241 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9728 N$19456 N$19455 "Straight Waveguide" sch_x=-241 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9729 N$19458 N$19457 "Straight Waveguide" sch_x=-241 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9730 N$19460 N$19459 "Straight Waveguide" sch_x=-241 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9731 N$19462 N$19461 "Straight Waveguide" sch_x=-241 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9732 N$19464 N$19463 "Straight Waveguide" sch_x=-241 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9733 N$19466 N$19465 "Straight Waveguide" sch_x=-241 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9734 N$19468 N$19467 "Straight Waveguide" sch_x=-241 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9735 N$19470 N$19469 "Straight Waveguide" sch_x=-241 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9736 N$19472 N$19471 "Straight Waveguide" sch_x=-241 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9737 N$19474 N$19473 "Straight Waveguide" sch_x=-241 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9738 N$19476 N$19475 "Straight Waveguide" sch_x=-241 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9739 N$19478 N$19477 "Straight Waveguide" sch_x=-241 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9740 N$19480 N$19479 "Straight Waveguide" sch_x=-241 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9741 N$19482 N$19481 "Straight Waveguide" sch_x=-241 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9742 N$19484 N$19483 "Straight Waveguide" sch_x=-241 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9743 N$19486 N$19485 "Straight Waveguide" sch_x=-241 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9744 N$19488 N$19487 "Straight Waveguide" sch_x=-241 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9745 N$19490 N$19489 "Straight Waveguide" sch_x=-241 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9746 N$19492 N$19491 "Straight Waveguide" sch_x=-241 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9747 N$19494 N$19493 "Straight Waveguide" sch_x=-241 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9748 N$19496 N$19495 "Straight Waveguide" sch_x=-241 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9749 N$19498 N$19497 "Straight Waveguide" sch_x=-241 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9750 N$19500 N$19499 "Straight Waveguide" sch_x=-241 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9751 N$19502 N$19501 "Straight Waveguide" sch_x=-241 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9752 N$19504 N$19503 "Straight Waveguide" sch_x=-241 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9753 N$19506 N$19505 "Straight Waveguide" sch_x=-241 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9754 N$19508 N$19507 "Straight Waveguide" sch_x=-241 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9755 N$19510 N$19509 "Straight Waveguide" sch_x=-241 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9756 N$19512 N$19511 "Straight Waveguide" sch_x=-241 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9757 N$19514 N$19513 "Straight Waveguide" sch_x=-241 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9758 N$19516 N$19515 "Straight Waveguide" sch_x=-241 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9759 N$19518 N$19517 "Straight Waveguide" sch_x=-241 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9760 N$19520 N$19519 "Straight Waveguide" sch_x=-241 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9761 N$19522 N$19521 "Straight Waveguide" sch_x=-241 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9762 N$19524 N$19523 "Straight Waveguide" sch_x=-241 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9763 N$19526 N$19525 "Straight Waveguide" sch_x=-241 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9764 N$19528 N$19527 "Straight Waveguide" sch_x=-241 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9765 N$19530 N$19529 "Straight Waveguide" sch_x=-241 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9766 N$19532 N$19531 "Straight Waveguide" sch_x=-241 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9767 N$19534 N$19533 "Straight Waveguide" sch_x=-241 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9768 N$19536 N$19535 "Straight Waveguide" sch_x=-241 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9769 N$19538 N$19537 "Straight Waveguide" sch_x=-241 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9770 N$19540 N$19539 "Straight Waveguide" sch_x=-241 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9771 N$19542 N$19541 "Straight Waveguide" sch_x=-241 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9772 N$19544 N$19543 "Straight Waveguide" sch_x=-241 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9773 N$19546 N$19545 "Straight Waveguide" sch_x=-241 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9774 N$19548 N$19547 "Straight Waveguide" sch_x=-241 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9775 N$19550 N$19549 "Straight Waveguide" sch_x=-241 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9776 N$19552 N$19551 "Straight Waveguide" sch_x=-241 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9777 N$19554 N$19553 "Straight Waveguide" sch_x=-241 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9778 N$19556 N$19555 "Straight Waveguide" sch_x=-241 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9779 N$19558 N$19557 "Straight Waveguide" sch_x=-241 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9780 N$19560 N$19559 "Straight Waveguide" sch_x=-241 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9781 N$19562 N$19561 "Straight Waveguide" sch_x=-241 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9782 N$19564 N$19563 "Straight Waveguide" sch_x=-241 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9783 N$19566 N$19565 "Straight Waveguide" sch_x=-241 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9784 N$19568 N$19567 "Straight Waveguide" sch_x=-241 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9785 N$19570 N$19569 "Straight Waveguide" sch_x=-241 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9786 N$19572 N$19571 "Straight Waveguide" sch_x=-241 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9787 N$19574 N$19573 "Straight Waveguide" sch_x=-241 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9788 N$19576 N$19575 "Straight Waveguide" sch_x=-241 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9789 N$19578 N$19577 "Straight Waveguide" sch_x=-241 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9790 N$19580 N$19579 "Straight Waveguide" sch_x=-241 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9791 N$19582 N$19581 "Straight Waveguide" sch_x=-241 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9792 N$19584 N$19583 "Straight Waveguide" sch_x=-241 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9793 N$19586 N$19585 "Straight Waveguide" sch_x=-241 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9794 N$19588 N$19587 "Straight Waveguide" sch_x=-241 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9795 N$19590 N$19589 "Straight Waveguide" sch_x=-241 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9796 N$19592 N$19591 "Straight Waveguide" sch_x=-241 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9797 N$19594 N$19593 "Straight Waveguide" sch_x=-241 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9798 N$19596 N$19595 "Straight Waveguide" sch_x=-241 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9799 N$19598 N$19597 "Straight Waveguide" sch_x=-241 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9800 N$19600 N$19599 "Straight Waveguide" sch_x=-241 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9801 N$19602 N$19601 "Straight Waveguide" sch_x=-239 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9802 N$19604 N$19603 "Straight Waveguide" sch_x=-239 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9803 N$19606 N$19605 "Straight Waveguide" sch_x=-239 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9804 N$19608 N$19607 "Straight Waveguide" sch_x=-239 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9805 N$19610 N$19609 "Straight Waveguide" sch_x=-239 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9806 N$19612 N$19611 "Straight Waveguide" sch_x=-239 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9807 N$19614 N$19613 "Straight Waveguide" sch_x=-239 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9808 N$19616 N$19615 "Straight Waveguide" sch_x=-239 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9809 N$19618 N$19617 "Straight Waveguide" sch_x=-239 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9810 N$19620 N$19619 "Straight Waveguide" sch_x=-239 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9811 N$19622 N$19621 "Straight Waveguide" sch_x=-239 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9812 N$19624 N$19623 "Straight Waveguide" sch_x=-239 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9813 N$19626 N$19625 "Straight Waveguide" sch_x=-239 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9814 N$19628 N$19627 "Straight Waveguide" sch_x=-239 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9815 N$19630 N$19629 "Straight Waveguide" sch_x=-239 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9816 N$19632 N$19631 "Straight Waveguide" sch_x=-239 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9817 N$19634 N$19633 "Straight Waveguide" sch_x=-239 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9818 N$19636 N$19635 "Straight Waveguide" sch_x=-239 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9819 N$19638 N$19637 "Straight Waveguide" sch_x=-239 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9820 N$19640 N$19639 "Straight Waveguide" sch_x=-239 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9821 N$19642 N$19641 "Straight Waveguide" sch_x=-239 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9822 N$19644 N$19643 "Straight Waveguide" sch_x=-239 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9823 N$19646 N$19645 "Straight Waveguide" sch_x=-239 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9824 N$19648 N$19647 "Straight Waveguide" sch_x=-239 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9825 N$19650 N$19649 "Straight Waveguide" sch_x=-239 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9826 N$19652 N$19651 "Straight Waveguide" sch_x=-239 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9827 N$19654 N$19653 "Straight Waveguide" sch_x=-239 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9828 N$19656 N$19655 "Straight Waveguide" sch_x=-239 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9829 N$19658 N$19657 "Straight Waveguide" sch_x=-239 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9830 N$19660 N$19659 "Straight Waveguide" sch_x=-239 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9831 N$19662 N$19661 "Straight Waveguide" sch_x=-239 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9832 N$19664 N$19663 "Straight Waveguide" sch_x=-239 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9833 N$19666 N$19665 "Straight Waveguide" sch_x=-239 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9834 N$19668 N$19667 "Straight Waveguide" sch_x=-239 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9835 N$19670 N$19669 "Straight Waveguide" sch_x=-239 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9836 N$19672 N$19671 "Straight Waveguide" sch_x=-239 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9837 N$19674 N$19673 "Straight Waveguide" sch_x=-239 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9838 N$19676 N$19675 "Straight Waveguide" sch_x=-239 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9839 N$19678 N$19677 "Straight Waveguide" sch_x=-239 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9840 N$19680 N$19679 "Straight Waveguide" sch_x=-239 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9841 N$19682 N$19681 "Straight Waveguide" sch_x=-239 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9842 N$19684 N$19683 "Straight Waveguide" sch_x=-239 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9843 N$19686 N$19685 "Straight Waveguide" sch_x=-239 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9844 N$19688 N$19687 "Straight Waveguide" sch_x=-239 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9845 N$19690 N$19689 "Straight Waveguide" sch_x=-239 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9846 N$19692 N$19691 "Straight Waveguide" sch_x=-239 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9847 N$19694 N$19693 "Straight Waveguide" sch_x=-239 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9848 N$19696 N$19695 "Straight Waveguide" sch_x=-239 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9849 N$19698 N$19697 "Straight Waveguide" sch_x=-239 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9850 N$19700 N$19699 "Straight Waveguide" sch_x=-239 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9851 N$19702 N$19701 "Straight Waveguide" sch_x=-239 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9852 N$19704 N$19703 "Straight Waveguide" sch_x=-239 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9853 N$19706 N$19705 "Straight Waveguide" sch_x=-239 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9854 N$19708 N$19707 "Straight Waveguide" sch_x=-239 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9855 N$19710 N$19709 "Straight Waveguide" sch_x=-239 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9856 N$19712 N$19711 "Straight Waveguide" sch_x=-239 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9857 N$19714 N$19713 "Straight Waveguide" sch_x=-239 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9858 N$19716 N$19715 "Straight Waveguide" sch_x=-239 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9859 N$19718 N$19717 "Straight Waveguide" sch_x=-239 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9860 N$19720 N$19719 "Straight Waveguide" sch_x=-239 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9861 N$19722 N$19721 "Straight Waveguide" sch_x=-239 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9862 N$19724 N$19723 "Straight Waveguide" sch_x=-239 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9863 N$19726 N$19725 "Straight Waveguide" sch_x=-239 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9864 N$19728 N$19727 "Straight Waveguide" sch_x=-239 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9865 N$19730 N$19729 "Straight Waveguide" sch_x=-239 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9866 N$19732 N$19731 "Straight Waveguide" sch_x=-239 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9867 N$19734 N$19733 "Straight Waveguide" sch_x=-239 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9868 N$19736 N$19735 "Straight Waveguide" sch_x=-239 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9869 N$19738 N$19737 "Straight Waveguide" sch_x=-239 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9870 N$19740 N$19739 "Straight Waveguide" sch_x=-239 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9871 N$19742 N$19741 "Straight Waveguide" sch_x=-239 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9872 N$19744 N$19743 "Straight Waveguide" sch_x=-239 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9873 N$19746 N$19745 "Straight Waveguide" sch_x=-239 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9874 N$19748 N$19747 "Straight Waveguide" sch_x=-239 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9875 N$19750 N$19749 "Straight Waveguide" sch_x=-239 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9876 N$19752 N$19751 "Straight Waveguide" sch_x=-239 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9877 N$19754 N$19753 "Straight Waveguide" sch_x=-239 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9878 N$19756 N$19755 "Straight Waveguide" sch_x=-239 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9879 N$19758 N$19757 "Straight Waveguide" sch_x=-239 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9880 N$19760 N$19759 "Straight Waveguide" sch_x=-239 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9881 N$19762 N$19761 "Straight Waveguide" sch_x=-239 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9882 N$19764 N$19763 "Straight Waveguide" sch_x=-239 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9883 N$19766 N$19765 "Straight Waveguide" sch_x=-239 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9884 N$19768 N$19767 "Straight Waveguide" sch_x=-239 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9885 N$19770 N$19769 "Straight Waveguide" sch_x=-239 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9886 N$19772 N$19771 "Straight Waveguide" sch_x=-239 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9887 N$19774 N$19773 "Straight Waveguide" sch_x=-239 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9888 N$19776 N$19775 "Straight Waveguide" sch_x=-239 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9889 N$19778 N$19777 "Straight Waveguide" sch_x=-239 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9890 N$19780 N$19779 "Straight Waveguide" sch_x=-239 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9891 N$19782 N$19781 "Straight Waveguide" sch_x=-239 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9892 N$19784 N$19783 "Straight Waveguide" sch_x=-239 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9893 N$19786 N$19785 "Straight Waveguide" sch_x=-239 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9894 N$19788 N$19787 "Straight Waveguide" sch_x=-239 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9895 N$19790 N$19789 "Straight Waveguide" sch_x=-239 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9896 N$19792 N$19791 "Straight Waveguide" sch_x=-239 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9897 N$19794 N$19793 "Straight Waveguide" sch_x=-239 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9898 N$19796 N$19795 "Straight Waveguide" sch_x=-239 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9899 N$19798 N$19797 "Straight Waveguide" sch_x=-239 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9900 N$19800 N$19799 "Straight Waveguide" sch_x=-239 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9901 N$19802 N$19801 "Straight Waveguide" sch_x=-239 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9902 N$19804 N$19803 "Straight Waveguide" sch_x=-239 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9903 N$19806 N$19805 "Straight Waveguide" sch_x=-239 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9904 N$19808 N$19807 "Straight Waveguide" sch_x=-239 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9905 N$19810 N$19809 "Straight Waveguide" sch_x=-239 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9906 N$19812 N$19811 "Straight Waveguide" sch_x=-239 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9907 N$19814 N$19813 "Straight Waveguide" sch_x=-239 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9908 N$19816 N$19815 "Straight Waveguide" sch_x=-239 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9909 N$19818 N$19817 "Straight Waveguide" sch_x=-239 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9910 N$19820 N$19819 "Straight Waveguide" sch_x=-239 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9911 N$19822 N$19821 "Straight Waveguide" sch_x=-239 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9912 N$19824 N$19823 "Straight Waveguide" sch_x=-239 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9913 N$19826 N$19825 "Straight Waveguide" sch_x=-237 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9914 N$19828 N$19827 "Straight Waveguide" sch_x=-237 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9915 N$19830 N$19829 "Straight Waveguide" sch_x=-237 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9916 N$19832 N$19831 "Straight Waveguide" sch_x=-237 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9917 N$19834 N$19833 "Straight Waveguide" sch_x=-237 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9918 N$19836 N$19835 "Straight Waveguide" sch_x=-237 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9919 N$19838 N$19837 "Straight Waveguide" sch_x=-237 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9920 N$19840 N$19839 "Straight Waveguide" sch_x=-237 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9921 N$19842 N$19841 "Straight Waveguide" sch_x=-237 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9922 N$19844 N$19843 "Straight Waveguide" sch_x=-237 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9923 N$19846 N$19845 "Straight Waveguide" sch_x=-237 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9924 N$19848 N$19847 "Straight Waveguide" sch_x=-237 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9925 N$19850 N$19849 "Straight Waveguide" sch_x=-237 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9926 N$19852 N$19851 "Straight Waveguide" sch_x=-237 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9927 N$19854 N$19853 "Straight Waveguide" sch_x=-237 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9928 N$19856 N$19855 "Straight Waveguide" sch_x=-237 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9929 N$19858 N$19857 "Straight Waveguide" sch_x=-237 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9930 N$19860 N$19859 "Straight Waveguide" sch_x=-237 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9931 N$19862 N$19861 "Straight Waveguide" sch_x=-237 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9932 N$19864 N$19863 "Straight Waveguide" sch_x=-237 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9933 N$19866 N$19865 "Straight Waveguide" sch_x=-237 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9934 N$19868 N$19867 "Straight Waveguide" sch_x=-237 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9935 N$19870 N$19869 "Straight Waveguide" sch_x=-237 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9936 N$19872 N$19871 "Straight Waveguide" sch_x=-237 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9937 N$19874 N$19873 "Straight Waveguide" sch_x=-237 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9938 N$19876 N$19875 "Straight Waveguide" sch_x=-237 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9939 N$19878 N$19877 "Straight Waveguide" sch_x=-237 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9940 N$19880 N$19879 "Straight Waveguide" sch_x=-237 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9941 N$19882 N$19881 "Straight Waveguide" sch_x=-237 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9942 N$19884 N$19883 "Straight Waveguide" sch_x=-237 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9943 N$19886 N$19885 "Straight Waveguide" sch_x=-237 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9944 N$19888 N$19887 "Straight Waveguide" sch_x=-237 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9945 N$19890 N$19889 "Straight Waveguide" sch_x=-237 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9946 N$19892 N$19891 "Straight Waveguide" sch_x=-237 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9947 N$19894 N$19893 "Straight Waveguide" sch_x=-237 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9948 N$19896 N$19895 "Straight Waveguide" sch_x=-237 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9949 N$19898 N$19897 "Straight Waveguide" sch_x=-237 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9950 N$19900 N$19899 "Straight Waveguide" sch_x=-237 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9951 N$19902 N$19901 "Straight Waveguide" sch_x=-237 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9952 N$19904 N$19903 "Straight Waveguide" sch_x=-237 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9953 N$19906 N$19905 "Straight Waveguide" sch_x=-237 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9954 N$19908 N$19907 "Straight Waveguide" sch_x=-237 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9955 N$19910 N$19909 "Straight Waveguide" sch_x=-237 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9956 N$19912 N$19911 "Straight Waveguide" sch_x=-237 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9957 N$19914 N$19913 "Straight Waveguide" sch_x=-237 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9958 N$19916 N$19915 "Straight Waveguide" sch_x=-237 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9959 N$19918 N$19917 "Straight Waveguide" sch_x=-237 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9960 N$19920 N$19919 "Straight Waveguide" sch_x=-237 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9961 N$19922 N$19921 "Straight Waveguide" sch_x=-237 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9962 N$19924 N$19923 "Straight Waveguide" sch_x=-237 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9963 N$19926 N$19925 "Straight Waveguide" sch_x=-237 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9964 N$19928 N$19927 "Straight Waveguide" sch_x=-237 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9965 N$19930 N$19929 "Straight Waveguide" sch_x=-237 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9966 N$19932 N$19931 "Straight Waveguide" sch_x=-237 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9967 N$19934 N$19933 "Straight Waveguide" sch_x=-237 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9968 N$19936 N$19935 "Straight Waveguide" sch_x=-237 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9969 N$19938 N$19937 "Straight Waveguide" sch_x=-237 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9970 N$19940 N$19939 "Straight Waveguide" sch_x=-237 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9971 N$19942 N$19941 "Straight Waveguide" sch_x=-237 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9972 N$19944 N$19943 "Straight Waveguide" sch_x=-237 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9973 N$19946 N$19945 "Straight Waveguide" sch_x=-237 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9974 N$19948 N$19947 "Straight Waveguide" sch_x=-237 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9975 N$19950 N$19949 "Straight Waveguide" sch_x=-237 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9976 N$19952 N$19951 "Straight Waveguide" sch_x=-237 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9977 N$19954 N$19953 "Straight Waveguide" sch_x=-237 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9978 N$19956 N$19955 "Straight Waveguide" sch_x=-237 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9979 N$19958 N$19957 "Straight Waveguide" sch_x=-237 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9980 N$19960 N$19959 "Straight Waveguide" sch_x=-237 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9981 N$19962 N$19961 "Straight Waveguide" sch_x=-237 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9982 N$19964 N$19963 "Straight Waveguide" sch_x=-237 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9983 N$19966 N$19965 "Straight Waveguide" sch_x=-237 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9984 N$19968 N$19967 "Straight Waveguide" sch_x=-237 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9985 N$19970 N$19969 "Straight Waveguide" sch_x=-237 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9986 N$19972 N$19971 "Straight Waveguide" sch_x=-237 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9987 N$19974 N$19973 "Straight Waveguide" sch_x=-237 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9988 N$19976 N$19975 "Straight Waveguide" sch_x=-237 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9989 N$19978 N$19977 "Straight Waveguide" sch_x=-237 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9990 N$19980 N$19979 "Straight Waveguide" sch_x=-237 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9991 N$19982 N$19981 "Straight Waveguide" sch_x=-237 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9992 N$19984 N$19983 "Straight Waveguide" sch_x=-237 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9993 N$19986 N$19985 "Straight Waveguide" sch_x=-237 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9994 N$19988 N$19987 "Straight Waveguide" sch_x=-237 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9995 N$19990 N$19989 "Straight Waveguide" sch_x=-237 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9996 N$19992 N$19991 "Straight Waveguide" sch_x=-237 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9997 N$19994 N$19993 "Straight Waveguide" sch_x=-237 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9998 N$19996 N$19995 "Straight Waveguide" sch_x=-237 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9999 N$19998 N$19997 "Straight Waveguide" sch_x=-237 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10000 N$20000 N$19999 "Straight Waveguide" sch_x=-237 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10001 N$20002 N$20001 "Straight Waveguide" sch_x=-237 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10002 N$20004 N$20003 "Straight Waveguide" sch_x=-237 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10003 N$20006 N$20005 "Straight Waveguide" sch_x=-237 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10004 N$20008 N$20007 "Straight Waveguide" sch_x=-237 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10005 N$20010 N$20009 "Straight Waveguide" sch_x=-237 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10006 N$20012 N$20011 "Straight Waveguide" sch_x=-237 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10007 N$20014 N$20013 "Straight Waveguide" sch_x=-237 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10008 N$20016 N$20015 "Straight Waveguide" sch_x=-237 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10009 N$20018 N$20017 "Straight Waveguide" sch_x=-237 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10010 N$20020 N$20019 "Straight Waveguide" sch_x=-237 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10011 N$20022 N$20021 "Straight Waveguide" sch_x=-237 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10012 N$20024 N$20023 "Straight Waveguide" sch_x=-237 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10013 N$20026 N$20025 "Straight Waveguide" sch_x=-237 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10014 N$20028 N$20027 "Straight Waveguide" sch_x=-237 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10015 N$20030 N$20029 "Straight Waveguide" sch_x=-237 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10016 N$20032 N$20031 "Straight Waveguide" sch_x=-237 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10017 N$20034 N$20033 "Straight Waveguide" sch_x=-237 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10018 N$20036 N$20035 "Straight Waveguide" sch_x=-237 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10019 N$20038 N$20037 "Straight Waveguide" sch_x=-237 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10020 N$20040 N$20039 "Straight Waveguide" sch_x=-237 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10021 N$20042 N$20041 "Straight Waveguide" sch_x=-237 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10022 N$20044 N$20043 "Straight Waveguide" sch_x=-237 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10023 N$20046 N$20045 "Straight Waveguide" sch_x=-235 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10024 N$20048 N$20047 "Straight Waveguide" sch_x=-235 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10025 N$20050 N$20049 "Straight Waveguide" sch_x=-235 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10026 N$20052 N$20051 "Straight Waveguide" sch_x=-235 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10027 N$20054 N$20053 "Straight Waveguide" sch_x=-235 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10028 N$20056 N$20055 "Straight Waveguide" sch_x=-235 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10029 N$20058 N$20057 "Straight Waveguide" sch_x=-235 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10030 N$20060 N$20059 "Straight Waveguide" sch_x=-235 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10031 N$20062 N$20061 "Straight Waveguide" sch_x=-235 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10032 N$20064 N$20063 "Straight Waveguide" sch_x=-235 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10033 N$20066 N$20065 "Straight Waveguide" sch_x=-235 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10034 N$20068 N$20067 "Straight Waveguide" sch_x=-235 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10035 N$20070 N$20069 "Straight Waveguide" sch_x=-235 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10036 N$20072 N$20071 "Straight Waveguide" sch_x=-235 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10037 N$20074 N$20073 "Straight Waveguide" sch_x=-235 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10038 N$20076 N$20075 "Straight Waveguide" sch_x=-235 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10039 N$20078 N$20077 "Straight Waveguide" sch_x=-235 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10040 N$20080 N$20079 "Straight Waveguide" sch_x=-235 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10041 N$20082 N$20081 "Straight Waveguide" sch_x=-235 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10042 N$20084 N$20083 "Straight Waveguide" sch_x=-235 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10043 N$20086 N$20085 "Straight Waveguide" sch_x=-235 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10044 N$20088 N$20087 "Straight Waveguide" sch_x=-235 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10045 N$20090 N$20089 "Straight Waveguide" sch_x=-235 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10046 N$20092 N$20091 "Straight Waveguide" sch_x=-235 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10047 N$20094 N$20093 "Straight Waveguide" sch_x=-235 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10048 N$20096 N$20095 "Straight Waveguide" sch_x=-235 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10049 N$20098 N$20097 "Straight Waveguide" sch_x=-235 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10050 N$20100 N$20099 "Straight Waveguide" sch_x=-235 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10051 N$20102 N$20101 "Straight Waveguide" sch_x=-235 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10052 N$20104 N$20103 "Straight Waveguide" sch_x=-235 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10053 N$20106 N$20105 "Straight Waveguide" sch_x=-235 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10054 N$20108 N$20107 "Straight Waveguide" sch_x=-235 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10055 N$20110 N$20109 "Straight Waveguide" sch_x=-235 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10056 N$20112 N$20111 "Straight Waveguide" sch_x=-235 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10057 N$20114 N$20113 "Straight Waveguide" sch_x=-235 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10058 N$20116 N$20115 "Straight Waveguide" sch_x=-235 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10059 N$20118 N$20117 "Straight Waveguide" sch_x=-235 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10060 N$20120 N$20119 "Straight Waveguide" sch_x=-235 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10061 N$20122 N$20121 "Straight Waveguide" sch_x=-235 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10062 N$20124 N$20123 "Straight Waveguide" sch_x=-235 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10063 N$20126 N$20125 "Straight Waveguide" sch_x=-235 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10064 N$20128 N$20127 "Straight Waveguide" sch_x=-235 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10065 N$20130 N$20129 "Straight Waveguide" sch_x=-235 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10066 N$20132 N$20131 "Straight Waveguide" sch_x=-235 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10067 N$20134 N$20133 "Straight Waveguide" sch_x=-235 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10068 N$20136 N$20135 "Straight Waveguide" sch_x=-235 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10069 N$20138 N$20137 "Straight Waveguide" sch_x=-235 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10070 N$20140 N$20139 "Straight Waveguide" sch_x=-235 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10071 N$20142 N$20141 "Straight Waveguide" sch_x=-235 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10072 N$20144 N$20143 "Straight Waveguide" sch_x=-235 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10073 N$20146 N$20145 "Straight Waveguide" sch_x=-235 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10074 N$20148 N$20147 "Straight Waveguide" sch_x=-235 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10075 N$20150 N$20149 "Straight Waveguide" sch_x=-235 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10076 N$20152 N$20151 "Straight Waveguide" sch_x=-235 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10077 N$20154 N$20153 "Straight Waveguide" sch_x=-235 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10078 N$20156 N$20155 "Straight Waveguide" sch_x=-235 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10079 N$20158 N$20157 "Straight Waveguide" sch_x=-235 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10080 N$20160 N$20159 "Straight Waveguide" sch_x=-235 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10081 N$20162 N$20161 "Straight Waveguide" sch_x=-235 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10082 N$20164 N$20163 "Straight Waveguide" sch_x=-235 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10083 N$20166 N$20165 "Straight Waveguide" sch_x=-235 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10084 N$20168 N$20167 "Straight Waveguide" sch_x=-235 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10085 N$20170 N$20169 "Straight Waveguide" sch_x=-235 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10086 N$20172 N$20171 "Straight Waveguide" sch_x=-235 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10087 N$20174 N$20173 "Straight Waveguide" sch_x=-235 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10088 N$20176 N$20175 "Straight Waveguide" sch_x=-235 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10089 N$20178 N$20177 "Straight Waveguide" sch_x=-235 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10090 N$20180 N$20179 "Straight Waveguide" sch_x=-235 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10091 N$20182 N$20181 "Straight Waveguide" sch_x=-235 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10092 N$20184 N$20183 "Straight Waveguide" sch_x=-235 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10093 N$20186 N$20185 "Straight Waveguide" sch_x=-235 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10094 N$20188 N$20187 "Straight Waveguide" sch_x=-235 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10095 N$20190 N$20189 "Straight Waveguide" sch_x=-235 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10096 N$20192 N$20191 "Straight Waveguide" sch_x=-235 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10097 N$20194 N$20193 "Straight Waveguide" sch_x=-235 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10098 N$20196 N$20195 "Straight Waveguide" sch_x=-235 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10099 N$20198 N$20197 "Straight Waveguide" sch_x=-235 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10100 N$20200 N$20199 "Straight Waveguide" sch_x=-235 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10101 N$20202 N$20201 "Straight Waveguide" sch_x=-235 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10102 N$20204 N$20203 "Straight Waveguide" sch_x=-235 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10103 N$20206 N$20205 "Straight Waveguide" sch_x=-235 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10104 N$20208 N$20207 "Straight Waveguide" sch_x=-235 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10105 N$20210 N$20209 "Straight Waveguide" sch_x=-235 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10106 N$20212 N$20211 "Straight Waveguide" sch_x=-235 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10107 N$20214 N$20213 "Straight Waveguide" sch_x=-235 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10108 N$20216 N$20215 "Straight Waveguide" sch_x=-235 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10109 N$20218 N$20217 "Straight Waveguide" sch_x=-235 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10110 N$20220 N$20219 "Straight Waveguide" sch_x=-235 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10111 N$20222 N$20221 "Straight Waveguide" sch_x=-235 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10112 N$20224 N$20223 "Straight Waveguide" sch_x=-235 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10113 N$20226 N$20225 "Straight Waveguide" sch_x=-235 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10114 N$20228 N$20227 "Straight Waveguide" sch_x=-235 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10115 N$20230 N$20229 "Straight Waveguide" sch_x=-235 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10116 N$20232 N$20231 "Straight Waveguide" sch_x=-235 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10117 N$20234 N$20233 "Straight Waveguide" sch_x=-235 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10118 N$20236 N$20235 "Straight Waveguide" sch_x=-235 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10119 N$20238 N$20237 "Straight Waveguide" sch_x=-235 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10120 N$20240 N$20239 "Straight Waveguide" sch_x=-235 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10121 N$20242 N$20241 "Straight Waveguide" sch_x=-235 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10122 N$20244 N$20243 "Straight Waveguide" sch_x=-235 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10123 N$20246 N$20245 "Straight Waveguide" sch_x=-235 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10124 N$20248 N$20247 "Straight Waveguide" sch_x=-235 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10125 N$20250 N$20249 "Straight Waveguide" sch_x=-235 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10126 N$20252 N$20251 "Straight Waveguide" sch_x=-235 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10127 N$20254 N$20253 "Straight Waveguide" sch_x=-235 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10128 N$20256 N$20255 "Straight Waveguide" sch_x=-235 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10129 N$20258 N$20257 "Straight Waveguide" sch_x=-235 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10130 N$20260 N$20259 "Straight Waveguide" sch_x=-235 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10131 N$20262 N$20261 "Straight Waveguide" sch_x=-233 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10132 N$20264 N$20263 "Straight Waveguide" sch_x=-233 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10133 N$20266 N$20265 "Straight Waveguide" sch_x=-233 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10134 N$20268 N$20267 "Straight Waveguide" sch_x=-233 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10135 N$20270 N$20269 "Straight Waveguide" sch_x=-233 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10136 N$20272 N$20271 "Straight Waveguide" sch_x=-233 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10137 N$20274 N$20273 "Straight Waveguide" sch_x=-233 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10138 N$20276 N$20275 "Straight Waveguide" sch_x=-233 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10139 N$20278 N$20277 "Straight Waveguide" sch_x=-233 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10140 N$20280 N$20279 "Straight Waveguide" sch_x=-233 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10141 N$20282 N$20281 "Straight Waveguide" sch_x=-233 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10142 N$20284 N$20283 "Straight Waveguide" sch_x=-233 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10143 N$20286 N$20285 "Straight Waveguide" sch_x=-233 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10144 N$20288 N$20287 "Straight Waveguide" sch_x=-233 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10145 N$20290 N$20289 "Straight Waveguide" sch_x=-233 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10146 N$20292 N$20291 "Straight Waveguide" sch_x=-233 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10147 N$20294 N$20293 "Straight Waveguide" sch_x=-233 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10148 N$20296 N$20295 "Straight Waveguide" sch_x=-233 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10149 N$20298 N$20297 "Straight Waveguide" sch_x=-233 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10150 N$20300 N$20299 "Straight Waveguide" sch_x=-233 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10151 N$20302 N$20301 "Straight Waveguide" sch_x=-233 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10152 N$20304 N$20303 "Straight Waveguide" sch_x=-233 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10153 N$20306 N$20305 "Straight Waveguide" sch_x=-233 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10154 N$20308 N$20307 "Straight Waveguide" sch_x=-233 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10155 N$20310 N$20309 "Straight Waveguide" sch_x=-233 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10156 N$20312 N$20311 "Straight Waveguide" sch_x=-233 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10157 N$20314 N$20313 "Straight Waveguide" sch_x=-233 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10158 N$20316 N$20315 "Straight Waveguide" sch_x=-233 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10159 N$20318 N$20317 "Straight Waveguide" sch_x=-233 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10160 N$20320 N$20319 "Straight Waveguide" sch_x=-233 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10161 N$20322 N$20321 "Straight Waveguide" sch_x=-233 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10162 N$20324 N$20323 "Straight Waveguide" sch_x=-233 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10163 N$20326 N$20325 "Straight Waveguide" sch_x=-233 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10164 N$20328 N$20327 "Straight Waveguide" sch_x=-233 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10165 N$20330 N$20329 "Straight Waveguide" sch_x=-233 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10166 N$20332 N$20331 "Straight Waveguide" sch_x=-233 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10167 N$20334 N$20333 "Straight Waveguide" sch_x=-233 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10168 N$20336 N$20335 "Straight Waveguide" sch_x=-233 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10169 N$20338 N$20337 "Straight Waveguide" sch_x=-233 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10170 N$20340 N$20339 "Straight Waveguide" sch_x=-233 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10171 N$20342 N$20341 "Straight Waveguide" sch_x=-233 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10172 N$20344 N$20343 "Straight Waveguide" sch_x=-233 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10173 N$20346 N$20345 "Straight Waveguide" sch_x=-233 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10174 N$20348 N$20347 "Straight Waveguide" sch_x=-233 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10175 N$20350 N$20349 "Straight Waveguide" sch_x=-233 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10176 N$20352 N$20351 "Straight Waveguide" sch_x=-233 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10177 N$20354 N$20353 "Straight Waveguide" sch_x=-233 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10178 N$20356 N$20355 "Straight Waveguide" sch_x=-233 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10179 N$20358 N$20357 "Straight Waveguide" sch_x=-233 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10180 N$20360 N$20359 "Straight Waveguide" sch_x=-233 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10181 N$20362 N$20361 "Straight Waveguide" sch_x=-233 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10182 N$20364 N$20363 "Straight Waveguide" sch_x=-233 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10183 N$20366 N$20365 "Straight Waveguide" sch_x=-233 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10184 N$20368 N$20367 "Straight Waveguide" sch_x=-233 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10185 N$20370 N$20369 "Straight Waveguide" sch_x=-233 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10186 N$20372 N$20371 "Straight Waveguide" sch_x=-233 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10187 N$20374 N$20373 "Straight Waveguide" sch_x=-233 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10188 N$20376 N$20375 "Straight Waveguide" sch_x=-233 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10189 N$20378 N$20377 "Straight Waveguide" sch_x=-233 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10190 N$20380 N$20379 "Straight Waveguide" sch_x=-233 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10191 N$20382 N$20381 "Straight Waveguide" sch_x=-233 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10192 N$20384 N$20383 "Straight Waveguide" sch_x=-233 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10193 N$20386 N$20385 "Straight Waveguide" sch_x=-233 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10194 N$20388 N$20387 "Straight Waveguide" sch_x=-233 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10195 N$20390 N$20389 "Straight Waveguide" sch_x=-233 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10196 N$20392 N$20391 "Straight Waveguide" sch_x=-233 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10197 N$20394 N$20393 "Straight Waveguide" sch_x=-233 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10198 N$20396 N$20395 "Straight Waveguide" sch_x=-233 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10199 N$20398 N$20397 "Straight Waveguide" sch_x=-233 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10200 N$20400 N$20399 "Straight Waveguide" sch_x=-233 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10201 N$20402 N$20401 "Straight Waveguide" sch_x=-233 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10202 N$20404 N$20403 "Straight Waveguide" sch_x=-233 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10203 N$20406 N$20405 "Straight Waveguide" sch_x=-233 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10204 N$20408 N$20407 "Straight Waveguide" sch_x=-233 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10205 N$20410 N$20409 "Straight Waveguide" sch_x=-233 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10206 N$20412 N$20411 "Straight Waveguide" sch_x=-233 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10207 N$20414 N$20413 "Straight Waveguide" sch_x=-233 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10208 N$20416 N$20415 "Straight Waveguide" sch_x=-233 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10209 N$20418 N$20417 "Straight Waveguide" sch_x=-233 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10210 N$20420 N$20419 "Straight Waveguide" sch_x=-233 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10211 N$20422 N$20421 "Straight Waveguide" sch_x=-233 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10212 N$20424 N$20423 "Straight Waveguide" sch_x=-233 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10213 N$20426 N$20425 "Straight Waveguide" sch_x=-233 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10214 N$20428 N$20427 "Straight Waveguide" sch_x=-233 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10215 N$20430 N$20429 "Straight Waveguide" sch_x=-233 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10216 N$20432 N$20431 "Straight Waveguide" sch_x=-233 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10217 N$20434 N$20433 "Straight Waveguide" sch_x=-233 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10218 N$20436 N$20435 "Straight Waveguide" sch_x=-233 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10219 N$20438 N$20437 "Straight Waveguide" sch_x=-233 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10220 N$20440 N$20439 "Straight Waveguide" sch_x=-233 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10221 N$20442 N$20441 "Straight Waveguide" sch_x=-233 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10222 N$20444 N$20443 "Straight Waveguide" sch_x=-233 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10223 N$20446 N$20445 "Straight Waveguide" sch_x=-233 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10224 N$20448 N$20447 "Straight Waveguide" sch_x=-233 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10225 N$20450 N$20449 "Straight Waveguide" sch_x=-233 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10226 N$20452 N$20451 "Straight Waveguide" sch_x=-233 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10227 N$20454 N$20453 "Straight Waveguide" sch_x=-233 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10228 N$20456 N$20455 "Straight Waveguide" sch_x=-233 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10229 N$20458 N$20457 "Straight Waveguide" sch_x=-233 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10230 N$20460 N$20459 "Straight Waveguide" sch_x=-233 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10231 N$20462 N$20461 "Straight Waveguide" sch_x=-233 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10232 N$20464 N$20463 "Straight Waveguide" sch_x=-233 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10233 N$20466 N$20465 "Straight Waveguide" sch_x=-233 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10234 N$20468 N$20467 "Straight Waveguide" sch_x=-233 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10235 N$20470 N$20469 "Straight Waveguide" sch_x=-233 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10236 N$20472 N$20471 "Straight Waveguide" sch_x=-233 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10237 N$20474 N$20473 "Straight Waveguide" sch_x=-231 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10238 N$20476 N$20475 "Straight Waveguide" sch_x=-231 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10239 N$20478 N$20477 "Straight Waveguide" sch_x=-231 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10240 N$20480 N$20479 "Straight Waveguide" sch_x=-231 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10241 N$20482 N$20481 "Straight Waveguide" sch_x=-231 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10242 N$20484 N$20483 "Straight Waveguide" sch_x=-231 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10243 N$20486 N$20485 "Straight Waveguide" sch_x=-231 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10244 N$20488 N$20487 "Straight Waveguide" sch_x=-231 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10245 N$20490 N$20489 "Straight Waveguide" sch_x=-231 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10246 N$20492 N$20491 "Straight Waveguide" sch_x=-231 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10247 N$20494 N$20493 "Straight Waveguide" sch_x=-231 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10248 N$20496 N$20495 "Straight Waveguide" sch_x=-231 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10249 N$20498 N$20497 "Straight Waveguide" sch_x=-231 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10250 N$20500 N$20499 "Straight Waveguide" sch_x=-231 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10251 N$20502 N$20501 "Straight Waveguide" sch_x=-231 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10252 N$20504 N$20503 "Straight Waveguide" sch_x=-231 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10253 N$20506 N$20505 "Straight Waveguide" sch_x=-231 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10254 N$20508 N$20507 "Straight Waveguide" sch_x=-231 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10255 N$20510 N$20509 "Straight Waveguide" sch_x=-231 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10256 N$20512 N$20511 "Straight Waveguide" sch_x=-231 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10257 N$20514 N$20513 "Straight Waveguide" sch_x=-231 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10258 N$20516 N$20515 "Straight Waveguide" sch_x=-231 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10259 N$20518 N$20517 "Straight Waveguide" sch_x=-231 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10260 N$20520 N$20519 "Straight Waveguide" sch_x=-231 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10261 N$20522 N$20521 "Straight Waveguide" sch_x=-231 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10262 N$20524 N$20523 "Straight Waveguide" sch_x=-231 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10263 N$20526 N$20525 "Straight Waveguide" sch_x=-231 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10264 N$20528 N$20527 "Straight Waveguide" sch_x=-231 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10265 N$20530 N$20529 "Straight Waveguide" sch_x=-231 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10266 N$20532 N$20531 "Straight Waveguide" sch_x=-231 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10267 N$20534 N$20533 "Straight Waveguide" sch_x=-231 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10268 N$20536 N$20535 "Straight Waveguide" sch_x=-231 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10269 N$20538 N$20537 "Straight Waveguide" sch_x=-231 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10270 N$20540 N$20539 "Straight Waveguide" sch_x=-231 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10271 N$20542 N$20541 "Straight Waveguide" sch_x=-231 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10272 N$20544 N$20543 "Straight Waveguide" sch_x=-231 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10273 N$20546 N$20545 "Straight Waveguide" sch_x=-231 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10274 N$20548 N$20547 "Straight Waveguide" sch_x=-231 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10275 N$20550 N$20549 "Straight Waveguide" sch_x=-231 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10276 N$20552 N$20551 "Straight Waveguide" sch_x=-231 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10277 N$20554 N$20553 "Straight Waveguide" sch_x=-231 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10278 N$20556 N$20555 "Straight Waveguide" sch_x=-231 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10279 N$20558 N$20557 "Straight Waveguide" sch_x=-231 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10280 N$20560 N$20559 "Straight Waveguide" sch_x=-231 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10281 N$20562 N$20561 "Straight Waveguide" sch_x=-231 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10282 N$20564 N$20563 "Straight Waveguide" sch_x=-231 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10283 N$20566 N$20565 "Straight Waveguide" sch_x=-231 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10284 N$20568 N$20567 "Straight Waveguide" sch_x=-231 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10285 N$20570 N$20569 "Straight Waveguide" sch_x=-231 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10286 N$20572 N$20571 "Straight Waveguide" sch_x=-231 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10287 N$20574 N$20573 "Straight Waveguide" sch_x=-231 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10288 N$20576 N$20575 "Straight Waveguide" sch_x=-231 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10289 N$20578 N$20577 "Straight Waveguide" sch_x=-231 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10290 N$20580 N$20579 "Straight Waveguide" sch_x=-231 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10291 N$20582 N$20581 "Straight Waveguide" sch_x=-231 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10292 N$20584 N$20583 "Straight Waveguide" sch_x=-231 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10293 N$20586 N$20585 "Straight Waveguide" sch_x=-231 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10294 N$20588 N$20587 "Straight Waveguide" sch_x=-231 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10295 N$20590 N$20589 "Straight Waveguide" sch_x=-231 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10296 N$20592 N$20591 "Straight Waveguide" sch_x=-231 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10297 N$20594 N$20593 "Straight Waveguide" sch_x=-231 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10298 N$20596 N$20595 "Straight Waveguide" sch_x=-231 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10299 N$20598 N$20597 "Straight Waveguide" sch_x=-231 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10300 N$20600 N$20599 "Straight Waveguide" sch_x=-231 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10301 N$20602 N$20601 "Straight Waveguide" sch_x=-231 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10302 N$20604 N$20603 "Straight Waveguide" sch_x=-231 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10303 N$20606 N$20605 "Straight Waveguide" sch_x=-231 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10304 N$20608 N$20607 "Straight Waveguide" sch_x=-231 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10305 N$20610 N$20609 "Straight Waveguide" sch_x=-231 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10306 N$20612 N$20611 "Straight Waveguide" sch_x=-231 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10307 N$20614 N$20613 "Straight Waveguide" sch_x=-231 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10308 N$20616 N$20615 "Straight Waveguide" sch_x=-231 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10309 N$20618 N$20617 "Straight Waveguide" sch_x=-231 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10310 N$20620 N$20619 "Straight Waveguide" sch_x=-231 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10311 N$20622 N$20621 "Straight Waveguide" sch_x=-231 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10312 N$20624 N$20623 "Straight Waveguide" sch_x=-231 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10313 N$20626 N$20625 "Straight Waveguide" sch_x=-231 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10314 N$20628 N$20627 "Straight Waveguide" sch_x=-231 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10315 N$20630 N$20629 "Straight Waveguide" sch_x=-231 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10316 N$20632 N$20631 "Straight Waveguide" sch_x=-231 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10317 N$20634 N$20633 "Straight Waveguide" sch_x=-231 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10318 N$20636 N$20635 "Straight Waveguide" sch_x=-231 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10319 N$20638 N$20637 "Straight Waveguide" sch_x=-231 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10320 N$20640 N$20639 "Straight Waveguide" sch_x=-231 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10321 N$20642 N$20641 "Straight Waveguide" sch_x=-231 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10322 N$20644 N$20643 "Straight Waveguide" sch_x=-231 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10323 N$20646 N$20645 "Straight Waveguide" sch_x=-231 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10324 N$20648 N$20647 "Straight Waveguide" sch_x=-231 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10325 N$20650 N$20649 "Straight Waveguide" sch_x=-231 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10326 N$20652 N$20651 "Straight Waveguide" sch_x=-231 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10327 N$20654 N$20653 "Straight Waveguide" sch_x=-231 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10328 N$20656 N$20655 "Straight Waveguide" sch_x=-231 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10329 N$20658 N$20657 "Straight Waveguide" sch_x=-231 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10330 N$20660 N$20659 "Straight Waveguide" sch_x=-231 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10331 N$20662 N$20661 "Straight Waveguide" sch_x=-231 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10332 N$20664 N$20663 "Straight Waveguide" sch_x=-231 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10333 N$20666 N$20665 "Straight Waveguide" sch_x=-231 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10334 N$20668 N$20667 "Straight Waveguide" sch_x=-231 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10335 N$20670 N$20669 "Straight Waveguide" sch_x=-231 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10336 N$20672 N$20671 "Straight Waveguide" sch_x=-231 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10337 N$20674 N$20673 "Straight Waveguide" sch_x=-231 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10338 N$20676 N$20675 "Straight Waveguide" sch_x=-231 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10339 N$20678 N$20677 "Straight Waveguide" sch_x=-231 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10340 N$20680 N$20679 "Straight Waveguide" sch_x=-231 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10341 N$20682 N$20681 "Straight Waveguide" sch_x=-229 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10342 N$20684 N$20683 "Straight Waveguide" sch_x=-229 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10343 N$20686 N$20685 "Straight Waveguide" sch_x=-229 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10344 N$20688 N$20687 "Straight Waveguide" sch_x=-229 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10345 N$20690 N$20689 "Straight Waveguide" sch_x=-229 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10346 N$20692 N$20691 "Straight Waveguide" sch_x=-229 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10347 N$20694 N$20693 "Straight Waveguide" sch_x=-229 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10348 N$20696 N$20695 "Straight Waveguide" sch_x=-229 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10349 N$20698 N$20697 "Straight Waveguide" sch_x=-229 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10350 N$20700 N$20699 "Straight Waveguide" sch_x=-229 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10351 N$20702 N$20701 "Straight Waveguide" sch_x=-229 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10352 N$20704 N$20703 "Straight Waveguide" sch_x=-229 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10353 N$20706 N$20705 "Straight Waveguide" sch_x=-229 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10354 N$20708 N$20707 "Straight Waveguide" sch_x=-229 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10355 N$20710 N$20709 "Straight Waveguide" sch_x=-229 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10356 N$20712 N$20711 "Straight Waveguide" sch_x=-229 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10357 N$20714 N$20713 "Straight Waveguide" sch_x=-229 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10358 N$20716 N$20715 "Straight Waveguide" sch_x=-229 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10359 N$20718 N$20717 "Straight Waveguide" sch_x=-229 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10360 N$20720 N$20719 "Straight Waveguide" sch_x=-229 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10361 N$20722 N$20721 "Straight Waveguide" sch_x=-229 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10362 N$20724 N$20723 "Straight Waveguide" sch_x=-229 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10363 N$20726 N$20725 "Straight Waveguide" sch_x=-229 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10364 N$20728 N$20727 "Straight Waveguide" sch_x=-229 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10365 N$20730 N$20729 "Straight Waveguide" sch_x=-229 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10366 N$20732 N$20731 "Straight Waveguide" sch_x=-229 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10367 N$20734 N$20733 "Straight Waveguide" sch_x=-229 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10368 N$20736 N$20735 "Straight Waveguide" sch_x=-229 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10369 N$20738 N$20737 "Straight Waveguide" sch_x=-229 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10370 N$20740 N$20739 "Straight Waveguide" sch_x=-229 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10371 N$20742 N$20741 "Straight Waveguide" sch_x=-229 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10372 N$20744 N$20743 "Straight Waveguide" sch_x=-229 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10373 N$20746 N$20745 "Straight Waveguide" sch_x=-229 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10374 N$20748 N$20747 "Straight Waveguide" sch_x=-229 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10375 N$20750 N$20749 "Straight Waveguide" sch_x=-229 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10376 N$20752 N$20751 "Straight Waveguide" sch_x=-229 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10377 N$20754 N$20753 "Straight Waveguide" sch_x=-229 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10378 N$20756 N$20755 "Straight Waveguide" sch_x=-229 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10379 N$20758 N$20757 "Straight Waveguide" sch_x=-229 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10380 N$20760 N$20759 "Straight Waveguide" sch_x=-229 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10381 N$20762 N$20761 "Straight Waveguide" sch_x=-229 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10382 N$20764 N$20763 "Straight Waveguide" sch_x=-229 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10383 N$20766 N$20765 "Straight Waveguide" sch_x=-229 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10384 N$20768 N$20767 "Straight Waveguide" sch_x=-229 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10385 N$20770 N$20769 "Straight Waveguide" sch_x=-229 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10386 N$20772 N$20771 "Straight Waveguide" sch_x=-229 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10387 N$20774 N$20773 "Straight Waveguide" sch_x=-229 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10388 N$20776 N$20775 "Straight Waveguide" sch_x=-229 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10389 N$20778 N$20777 "Straight Waveguide" sch_x=-229 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10390 N$20780 N$20779 "Straight Waveguide" sch_x=-229 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10391 N$20782 N$20781 "Straight Waveguide" sch_x=-229 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10392 N$20784 N$20783 "Straight Waveguide" sch_x=-229 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10393 N$20786 N$20785 "Straight Waveguide" sch_x=-229 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10394 N$20788 N$20787 "Straight Waveguide" sch_x=-229 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10395 N$20790 N$20789 "Straight Waveguide" sch_x=-229 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10396 N$20792 N$20791 "Straight Waveguide" sch_x=-229 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10397 N$20794 N$20793 "Straight Waveguide" sch_x=-229 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10398 N$20796 N$20795 "Straight Waveguide" sch_x=-229 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10399 N$20798 N$20797 "Straight Waveguide" sch_x=-229 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10400 N$20800 N$20799 "Straight Waveguide" sch_x=-229 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10401 N$20802 N$20801 "Straight Waveguide" sch_x=-229 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10402 N$20804 N$20803 "Straight Waveguide" sch_x=-229 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10403 N$20806 N$20805 "Straight Waveguide" sch_x=-229 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10404 N$20808 N$20807 "Straight Waveguide" sch_x=-229 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10405 N$20810 N$20809 "Straight Waveguide" sch_x=-229 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10406 N$20812 N$20811 "Straight Waveguide" sch_x=-229 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10407 N$20814 N$20813 "Straight Waveguide" sch_x=-229 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10408 N$20816 N$20815 "Straight Waveguide" sch_x=-229 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10409 N$20818 N$20817 "Straight Waveguide" sch_x=-229 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10410 N$20820 N$20819 "Straight Waveguide" sch_x=-229 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10411 N$20822 N$20821 "Straight Waveguide" sch_x=-229 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10412 N$20824 N$20823 "Straight Waveguide" sch_x=-229 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10413 N$20826 N$20825 "Straight Waveguide" sch_x=-229 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10414 N$20828 N$20827 "Straight Waveguide" sch_x=-229 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10415 N$20830 N$20829 "Straight Waveguide" sch_x=-229 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10416 N$20832 N$20831 "Straight Waveguide" sch_x=-229 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10417 N$20834 N$20833 "Straight Waveguide" sch_x=-229 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10418 N$20836 N$20835 "Straight Waveguide" sch_x=-229 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10419 N$20838 N$20837 "Straight Waveguide" sch_x=-229 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10420 N$20840 N$20839 "Straight Waveguide" sch_x=-229 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10421 N$20842 N$20841 "Straight Waveguide" sch_x=-229 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10422 N$20844 N$20843 "Straight Waveguide" sch_x=-229 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10423 N$20846 N$20845 "Straight Waveguide" sch_x=-229 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10424 N$20848 N$20847 "Straight Waveguide" sch_x=-229 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10425 N$20850 N$20849 "Straight Waveguide" sch_x=-229 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10426 N$20852 N$20851 "Straight Waveguide" sch_x=-229 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10427 N$20854 N$20853 "Straight Waveguide" sch_x=-229 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10428 N$20856 N$20855 "Straight Waveguide" sch_x=-229 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10429 N$20858 N$20857 "Straight Waveguide" sch_x=-229 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10430 N$20860 N$20859 "Straight Waveguide" sch_x=-229 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10431 N$20862 N$20861 "Straight Waveguide" sch_x=-229 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10432 N$20864 N$20863 "Straight Waveguide" sch_x=-229 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10433 N$20866 N$20865 "Straight Waveguide" sch_x=-229 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10434 N$20868 N$20867 "Straight Waveguide" sch_x=-229 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10435 N$20870 N$20869 "Straight Waveguide" sch_x=-229 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10436 N$20872 N$20871 "Straight Waveguide" sch_x=-229 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10437 N$20874 N$20873 "Straight Waveguide" sch_x=-229 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10438 N$20876 N$20875 "Straight Waveguide" sch_x=-229 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10439 N$20878 N$20877 "Straight Waveguide" sch_x=-229 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10440 N$20880 N$20879 "Straight Waveguide" sch_x=-229 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10441 N$20882 N$20881 "Straight Waveguide" sch_x=-229 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10442 N$20884 N$20883 "Straight Waveguide" sch_x=-229 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10443 N$20886 N$20885 "Straight Waveguide" sch_x=-227 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10444 N$20888 N$20887 "Straight Waveguide" sch_x=-227 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10445 N$20890 N$20889 "Straight Waveguide" sch_x=-227 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10446 N$20892 N$20891 "Straight Waveguide" sch_x=-227 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10447 N$20894 N$20893 "Straight Waveguide" sch_x=-227 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10448 N$20896 N$20895 "Straight Waveguide" sch_x=-227 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10449 N$20898 N$20897 "Straight Waveguide" sch_x=-227 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10450 N$20900 N$20899 "Straight Waveguide" sch_x=-227 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10451 N$20902 N$20901 "Straight Waveguide" sch_x=-227 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10452 N$20904 N$20903 "Straight Waveguide" sch_x=-227 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10453 N$20906 N$20905 "Straight Waveguide" sch_x=-227 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10454 N$20908 N$20907 "Straight Waveguide" sch_x=-227 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10455 N$20910 N$20909 "Straight Waveguide" sch_x=-227 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10456 N$20912 N$20911 "Straight Waveguide" sch_x=-227 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10457 N$20914 N$20913 "Straight Waveguide" sch_x=-227 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10458 N$20916 N$20915 "Straight Waveguide" sch_x=-227 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10459 N$20918 N$20917 "Straight Waveguide" sch_x=-227 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10460 N$20920 N$20919 "Straight Waveguide" sch_x=-227 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10461 N$20922 N$20921 "Straight Waveguide" sch_x=-227 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10462 N$20924 N$20923 "Straight Waveguide" sch_x=-227 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10463 N$20926 N$20925 "Straight Waveguide" sch_x=-227 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10464 N$20928 N$20927 "Straight Waveguide" sch_x=-227 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10465 N$20930 N$20929 "Straight Waveguide" sch_x=-227 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10466 N$20932 N$20931 "Straight Waveguide" sch_x=-227 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10467 N$20934 N$20933 "Straight Waveguide" sch_x=-227 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10468 N$20936 N$20935 "Straight Waveguide" sch_x=-227 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10469 N$20938 N$20937 "Straight Waveguide" sch_x=-227 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10470 N$20940 N$20939 "Straight Waveguide" sch_x=-227 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10471 N$20942 N$20941 "Straight Waveguide" sch_x=-227 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10472 N$20944 N$20943 "Straight Waveguide" sch_x=-227 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10473 N$20946 N$20945 "Straight Waveguide" sch_x=-227 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10474 N$20948 N$20947 "Straight Waveguide" sch_x=-227 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10475 N$20950 N$20949 "Straight Waveguide" sch_x=-227 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10476 N$20952 N$20951 "Straight Waveguide" sch_x=-227 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10477 N$20954 N$20953 "Straight Waveguide" sch_x=-227 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10478 N$20956 N$20955 "Straight Waveguide" sch_x=-227 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10479 N$20958 N$20957 "Straight Waveguide" sch_x=-227 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10480 N$20960 N$20959 "Straight Waveguide" sch_x=-227 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10481 N$20962 N$20961 "Straight Waveguide" sch_x=-227 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10482 N$20964 N$20963 "Straight Waveguide" sch_x=-227 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10483 N$20966 N$20965 "Straight Waveguide" sch_x=-227 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10484 N$20968 N$20967 "Straight Waveguide" sch_x=-227 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10485 N$20970 N$20969 "Straight Waveguide" sch_x=-227 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10486 N$20972 N$20971 "Straight Waveguide" sch_x=-227 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10487 N$20974 N$20973 "Straight Waveguide" sch_x=-227 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10488 N$20976 N$20975 "Straight Waveguide" sch_x=-227 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10489 N$20978 N$20977 "Straight Waveguide" sch_x=-227 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10490 N$20980 N$20979 "Straight Waveguide" sch_x=-227 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10491 N$20982 N$20981 "Straight Waveguide" sch_x=-227 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10492 N$20984 N$20983 "Straight Waveguide" sch_x=-227 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10493 N$20986 N$20985 "Straight Waveguide" sch_x=-227 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10494 N$20988 N$20987 "Straight Waveguide" sch_x=-227 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10495 N$20990 N$20989 "Straight Waveguide" sch_x=-227 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10496 N$20992 N$20991 "Straight Waveguide" sch_x=-227 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10497 N$20994 N$20993 "Straight Waveguide" sch_x=-227 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10498 N$20996 N$20995 "Straight Waveguide" sch_x=-227 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10499 N$20998 N$20997 "Straight Waveguide" sch_x=-227 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10500 N$21000 N$20999 "Straight Waveguide" sch_x=-227 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10501 N$21002 N$21001 "Straight Waveguide" sch_x=-227 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10502 N$21004 N$21003 "Straight Waveguide" sch_x=-227 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10503 N$21006 N$21005 "Straight Waveguide" sch_x=-227 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10504 N$21008 N$21007 "Straight Waveguide" sch_x=-227 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10505 N$21010 N$21009 "Straight Waveguide" sch_x=-227 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10506 N$21012 N$21011 "Straight Waveguide" sch_x=-227 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10507 N$21014 N$21013 "Straight Waveguide" sch_x=-227 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10508 N$21016 N$21015 "Straight Waveguide" sch_x=-227 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10509 N$21018 N$21017 "Straight Waveguide" sch_x=-227 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10510 N$21020 N$21019 "Straight Waveguide" sch_x=-227 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10511 N$21022 N$21021 "Straight Waveguide" sch_x=-227 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10512 N$21024 N$21023 "Straight Waveguide" sch_x=-227 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10513 N$21026 N$21025 "Straight Waveguide" sch_x=-227 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10514 N$21028 N$21027 "Straight Waveguide" sch_x=-227 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10515 N$21030 N$21029 "Straight Waveguide" sch_x=-227 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10516 N$21032 N$21031 "Straight Waveguide" sch_x=-227 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10517 N$21034 N$21033 "Straight Waveguide" sch_x=-227 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10518 N$21036 N$21035 "Straight Waveguide" sch_x=-227 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10519 N$21038 N$21037 "Straight Waveguide" sch_x=-227 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10520 N$21040 N$21039 "Straight Waveguide" sch_x=-227 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10521 N$21042 N$21041 "Straight Waveguide" sch_x=-227 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10522 N$21044 N$21043 "Straight Waveguide" sch_x=-227 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10523 N$21046 N$21045 "Straight Waveguide" sch_x=-227 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10524 N$21048 N$21047 "Straight Waveguide" sch_x=-227 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10525 N$21050 N$21049 "Straight Waveguide" sch_x=-227 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10526 N$21052 N$21051 "Straight Waveguide" sch_x=-227 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10527 N$21054 N$21053 "Straight Waveguide" sch_x=-227 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10528 N$21056 N$21055 "Straight Waveguide" sch_x=-227 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10529 N$21058 N$21057 "Straight Waveguide" sch_x=-227 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10530 N$21060 N$21059 "Straight Waveguide" sch_x=-227 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10531 N$21062 N$21061 "Straight Waveguide" sch_x=-227 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10532 N$21064 N$21063 "Straight Waveguide" sch_x=-227 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10533 N$21066 N$21065 "Straight Waveguide" sch_x=-227 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10534 N$21068 N$21067 "Straight Waveguide" sch_x=-227 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10535 N$21070 N$21069 "Straight Waveguide" sch_x=-227 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10536 N$21072 N$21071 "Straight Waveguide" sch_x=-227 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10537 N$21074 N$21073 "Straight Waveguide" sch_x=-227 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10538 N$21076 N$21075 "Straight Waveguide" sch_x=-227 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10539 N$21078 N$21077 "Straight Waveguide" sch_x=-227 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10540 N$21080 N$21079 "Straight Waveguide" sch_x=-227 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10541 N$21082 N$21081 "Straight Waveguide" sch_x=-227 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10542 N$21084 N$21083 "Straight Waveguide" sch_x=-227 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10543 N$21086 N$21085 "Straight Waveguide" sch_x=-225 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10544 N$21088 N$21087 "Straight Waveguide" sch_x=-225 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10545 N$21090 N$21089 "Straight Waveguide" sch_x=-225 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10546 N$21092 N$21091 "Straight Waveguide" sch_x=-225 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10547 N$21094 N$21093 "Straight Waveguide" sch_x=-225 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10548 N$21096 N$21095 "Straight Waveguide" sch_x=-225 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10549 N$21098 N$21097 "Straight Waveguide" sch_x=-225 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10550 N$21100 N$21099 "Straight Waveguide" sch_x=-225 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10551 N$21102 N$21101 "Straight Waveguide" sch_x=-225 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10552 N$21104 N$21103 "Straight Waveguide" sch_x=-225 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10553 N$21106 N$21105 "Straight Waveguide" sch_x=-225 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10554 N$21108 N$21107 "Straight Waveguide" sch_x=-225 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10555 N$21110 N$21109 "Straight Waveguide" sch_x=-225 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10556 N$21112 N$21111 "Straight Waveguide" sch_x=-225 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10557 N$21114 N$21113 "Straight Waveguide" sch_x=-225 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10558 N$21116 N$21115 "Straight Waveguide" sch_x=-225 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10559 N$21118 N$21117 "Straight Waveguide" sch_x=-225 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10560 N$21120 N$21119 "Straight Waveguide" sch_x=-225 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10561 N$21122 N$21121 "Straight Waveguide" sch_x=-225 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10562 N$21124 N$21123 "Straight Waveguide" sch_x=-225 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10563 N$21126 N$21125 "Straight Waveguide" sch_x=-225 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10564 N$21128 N$21127 "Straight Waveguide" sch_x=-225 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10565 N$21130 N$21129 "Straight Waveguide" sch_x=-225 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10566 N$21132 N$21131 "Straight Waveguide" sch_x=-225 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10567 N$21134 N$21133 "Straight Waveguide" sch_x=-225 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10568 N$21136 N$21135 "Straight Waveguide" sch_x=-225 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10569 N$21138 N$21137 "Straight Waveguide" sch_x=-225 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10570 N$21140 N$21139 "Straight Waveguide" sch_x=-225 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10571 N$21142 N$21141 "Straight Waveguide" sch_x=-225 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10572 N$21144 N$21143 "Straight Waveguide" sch_x=-225 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10573 N$21146 N$21145 "Straight Waveguide" sch_x=-225 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10574 N$21148 N$21147 "Straight Waveguide" sch_x=-225 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10575 N$21150 N$21149 "Straight Waveguide" sch_x=-225 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10576 N$21152 N$21151 "Straight Waveguide" sch_x=-225 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10577 N$21154 N$21153 "Straight Waveguide" sch_x=-225 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10578 N$21156 N$21155 "Straight Waveguide" sch_x=-225 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10579 N$21158 N$21157 "Straight Waveguide" sch_x=-225 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10580 N$21160 N$21159 "Straight Waveguide" sch_x=-225 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10581 N$21162 N$21161 "Straight Waveguide" sch_x=-225 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10582 N$21164 N$21163 "Straight Waveguide" sch_x=-225 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10583 N$21166 N$21165 "Straight Waveguide" sch_x=-225 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10584 N$21168 N$21167 "Straight Waveguide" sch_x=-225 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10585 N$21170 N$21169 "Straight Waveguide" sch_x=-225 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10586 N$21172 N$21171 "Straight Waveguide" sch_x=-225 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10587 N$21174 N$21173 "Straight Waveguide" sch_x=-225 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10588 N$21176 N$21175 "Straight Waveguide" sch_x=-225 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10589 N$21178 N$21177 "Straight Waveguide" sch_x=-225 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10590 N$21180 N$21179 "Straight Waveguide" sch_x=-225 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10591 N$21182 N$21181 "Straight Waveguide" sch_x=-225 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10592 N$21184 N$21183 "Straight Waveguide" sch_x=-225 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10593 N$21186 N$21185 "Straight Waveguide" sch_x=-225 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10594 N$21188 N$21187 "Straight Waveguide" sch_x=-225 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10595 N$21190 N$21189 "Straight Waveguide" sch_x=-225 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10596 N$21192 N$21191 "Straight Waveguide" sch_x=-225 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10597 N$21194 N$21193 "Straight Waveguide" sch_x=-225 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10598 N$21196 N$21195 "Straight Waveguide" sch_x=-225 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10599 N$21198 N$21197 "Straight Waveguide" sch_x=-225 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10600 N$21200 N$21199 "Straight Waveguide" sch_x=-225 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10601 N$21202 N$21201 "Straight Waveguide" sch_x=-225 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10602 N$21204 N$21203 "Straight Waveguide" sch_x=-225 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10603 N$21206 N$21205 "Straight Waveguide" sch_x=-225 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10604 N$21208 N$21207 "Straight Waveguide" sch_x=-225 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10605 N$21210 N$21209 "Straight Waveguide" sch_x=-225 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10606 N$21212 N$21211 "Straight Waveguide" sch_x=-225 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10607 N$21214 N$21213 "Straight Waveguide" sch_x=-225 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10608 N$21216 N$21215 "Straight Waveguide" sch_x=-225 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10609 N$21218 N$21217 "Straight Waveguide" sch_x=-225 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10610 N$21220 N$21219 "Straight Waveguide" sch_x=-225 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10611 N$21222 N$21221 "Straight Waveguide" sch_x=-225 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10612 N$21224 N$21223 "Straight Waveguide" sch_x=-225 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10613 N$21226 N$21225 "Straight Waveguide" sch_x=-225 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10614 N$21228 N$21227 "Straight Waveguide" sch_x=-225 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10615 N$21230 N$21229 "Straight Waveguide" sch_x=-225 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10616 N$21232 N$21231 "Straight Waveguide" sch_x=-225 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10617 N$21234 N$21233 "Straight Waveguide" sch_x=-225 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10618 N$21236 N$21235 "Straight Waveguide" sch_x=-225 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10619 N$21238 N$21237 "Straight Waveguide" sch_x=-225 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10620 N$21240 N$21239 "Straight Waveguide" sch_x=-225 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10621 N$21242 N$21241 "Straight Waveguide" sch_x=-225 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10622 N$21244 N$21243 "Straight Waveguide" sch_x=-225 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10623 N$21246 N$21245 "Straight Waveguide" sch_x=-225 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10624 N$21248 N$21247 "Straight Waveguide" sch_x=-225 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10625 N$21250 N$21249 "Straight Waveguide" sch_x=-225 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10626 N$21252 N$21251 "Straight Waveguide" sch_x=-225 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10627 N$21254 N$21253 "Straight Waveguide" sch_x=-225 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10628 N$21256 N$21255 "Straight Waveguide" sch_x=-225 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10629 N$21258 N$21257 "Straight Waveguide" sch_x=-225 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10630 N$21260 N$21259 "Straight Waveguide" sch_x=-225 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10631 N$21262 N$21261 "Straight Waveguide" sch_x=-225 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10632 N$21264 N$21263 "Straight Waveguide" sch_x=-225 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10633 N$21266 N$21265 "Straight Waveguide" sch_x=-225 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10634 N$21268 N$21267 "Straight Waveguide" sch_x=-225 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10635 N$21270 N$21269 "Straight Waveguide" sch_x=-225 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10636 N$21272 N$21271 "Straight Waveguide" sch_x=-225 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10637 N$21274 N$21273 "Straight Waveguide" sch_x=-225 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10638 N$21276 N$21275 "Straight Waveguide" sch_x=-225 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10639 N$21278 N$21277 "Straight Waveguide" sch_x=-225 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10640 N$21280 N$21279 "Straight Waveguide" sch_x=-225 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10641 N$21282 N$21281 "Straight Waveguide" sch_x=-223 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10642 N$21284 N$21283 "Straight Waveguide" sch_x=-223 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10643 N$21286 N$21285 "Straight Waveguide" sch_x=-223 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10644 N$21288 N$21287 "Straight Waveguide" sch_x=-223 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10645 N$21290 N$21289 "Straight Waveguide" sch_x=-223 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10646 N$21292 N$21291 "Straight Waveguide" sch_x=-223 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10647 N$21294 N$21293 "Straight Waveguide" sch_x=-223 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10648 N$21296 N$21295 "Straight Waveguide" sch_x=-223 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10649 N$21298 N$21297 "Straight Waveguide" sch_x=-223 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10650 N$21300 N$21299 "Straight Waveguide" sch_x=-223 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10651 N$21302 N$21301 "Straight Waveguide" sch_x=-223 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10652 N$21304 N$21303 "Straight Waveguide" sch_x=-223 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10653 N$21306 N$21305 "Straight Waveguide" sch_x=-223 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10654 N$21308 N$21307 "Straight Waveguide" sch_x=-223 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10655 N$21310 N$21309 "Straight Waveguide" sch_x=-223 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10656 N$21312 N$21311 "Straight Waveguide" sch_x=-223 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10657 N$21314 N$21313 "Straight Waveguide" sch_x=-223 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10658 N$21316 N$21315 "Straight Waveguide" sch_x=-223 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10659 N$21318 N$21317 "Straight Waveguide" sch_x=-223 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10660 N$21320 N$21319 "Straight Waveguide" sch_x=-223 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10661 N$21322 N$21321 "Straight Waveguide" sch_x=-223 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10662 N$21324 N$21323 "Straight Waveguide" sch_x=-223 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10663 N$21326 N$21325 "Straight Waveguide" sch_x=-223 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10664 N$21328 N$21327 "Straight Waveguide" sch_x=-223 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10665 N$21330 N$21329 "Straight Waveguide" sch_x=-223 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10666 N$21332 N$21331 "Straight Waveguide" sch_x=-223 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10667 N$21334 N$21333 "Straight Waveguide" sch_x=-223 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10668 N$21336 N$21335 "Straight Waveguide" sch_x=-223 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10669 N$21338 N$21337 "Straight Waveguide" sch_x=-223 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10670 N$21340 N$21339 "Straight Waveguide" sch_x=-223 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10671 N$21342 N$21341 "Straight Waveguide" sch_x=-223 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10672 N$21344 N$21343 "Straight Waveguide" sch_x=-223 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10673 N$21346 N$21345 "Straight Waveguide" sch_x=-223 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10674 N$21348 N$21347 "Straight Waveguide" sch_x=-223 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10675 N$21350 N$21349 "Straight Waveguide" sch_x=-223 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10676 N$21352 N$21351 "Straight Waveguide" sch_x=-223 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10677 N$21354 N$21353 "Straight Waveguide" sch_x=-223 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10678 N$21356 N$21355 "Straight Waveguide" sch_x=-223 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10679 N$21358 N$21357 "Straight Waveguide" sch_x=-223 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10680 N$21360 N$21359 "Straight Waveguide" sch_x=-223 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10681 N$21362 N$21361 "Straight Waveguide" sch_x=-223 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10682 N$21364 N$21363 "Straight Waveguide" sch_x=-223 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10683 N$21366 N$21365 "Straight Waveguide" sch_x=-223 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10684 N$21368 N$21367 "Straight Waveguide" sch_x=-223 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10685 N$21370 N$21369 "Straight Waveguide" sch_x=-223 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10686 N$21372 N$21371 "Straight Waveguide" sch_x=-223 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10687 N$21374 N$21373 "Straight Waveguide" sch_x=-223 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10688 N$21376 N$21375 "Straight Waveguide" sch_x=-223 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10689 N$21378 N$21377 "Straight Waveguide" sch_x=-223 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10690 N$21380 N$21379 "Straight Waveguide" sch_x=-223 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10691 N$21382 N$21381 "Straight Waveguide" sch_x=-223 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10692 N$21384 N$21383 "Straight Waveguide" sch_x=-223 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10693 N$21386 N$21385 "Straight Waveguide" sch_x=-223 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10694 N$21388 N$21387 "Straight Waveguide" sch_x=-223 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10695 N$21390 N$21389 "Straight Waveguide" sch_x=-223 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10696 N$21392 N$21391 "Straight Waveguide" sch_x=-223 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10697 N$21394 N$21393 "Straight Waveguide" sch_x=-223 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10698 N$21396 N$21395 "Straight Waveguide" sch_x=-223 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10699 N$21398 N$21397 "Straight Waveguide" sch_x=-223 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10700 N$21400 N$21399 "Straight Waveguide" sch_x=-223 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10701 N$21402 N$21401 "Straight Waveguide" sch_x=-223 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10702 N$21404 N$21403 "Straight Waveguide" sch_x=-223 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10703 N$21406 N$21405 "Straight Waveguide" sch_x=-223 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10704 N$21408 N$21407 "Straight Waveguide" sch_x=-223 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10705 N$21410 N$21409 "Straight Waveguide" sch_x=-223 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10706 N$21412 N$21411 "Straight Waveguide" sch_x=-223 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10707 N$21414 N$21413 "Straight Waveguide" sch_x=-223 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10708 N$21416 N$21415 "Straight Waveguide" sch_x=-223 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10709 N$21418 N$21417 "Straight Waveguide" sch_x=-223 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10710 N$21420 N$21419 "Straight Waveguide" sch_x=-223 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10711 N$21422 N$21421 "Straight Waveguide" sch_x=-223 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10712 N$21424 N$21423 "Straight Waveguide" sch_x=-223 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10713 N$21426 N$21425 "Straight Waveguide" sch_x=-223 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10714 N$21428 N$21427 "Straight Waveguide" sch_x=-223 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10715 N$21430 N$21429 "Straight Waveguide" sch_x=-223 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10716 N$21432 N$21431 "Straight Waveguide" sch_x=-223 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10717 N$21434 N$21433 "Straight Waveguide" sch_x=-223 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10718 N$21436 N$21435 "Straight Waveguide" sch_x=-223 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10719 N$21438 N$21437 "Straight Waveguide" sch_x=-223 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10720 N$21440 N$21439 "Straight Waveguide" sch_x=-223 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10721 N$21442 N$21441 "Straight Waveguide" sch_x=-223 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10722 N$21444 N$21443 "Straight Waveguide" sch_x=-223 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10723 N$21446 N$21445 "Straight Waveguide" sch_x=-223 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10724 N$21448 N$21447 "Straight Waveguide" sch_x=-223 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10725 N$21450 N$21449 "Straight Waveguide" sch_x=-223 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10726 N$21452 N$21451 "Straight Waveguide" sch_x=-223 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10727 N$21454 N$21453 "Straight Waveguide" sch_x=-223 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10728 N$21456 N$21455 "Straight Waveguide" sch_x=-223 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10729 N$21458 N$21457 "Straight Waveguide" sch_x=-223 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10730 N$21460 N$21459 "Straight Waveguide" sch_x=-223 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10731 N$21462 N$21461 "Straight Waveguide" sch_x=-223 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10732 N$21464 N$21463 "Straight Waveguide" sch_x=-223 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10733 N$21466 N$21465 "Straight Waveguide" sch_x=-223 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10734 N$21468 N$21467 "Straight Waveguide" sch_x=-223 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10735 N$21470 N$21469 "Straight Waveguide" sch_x=-223 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10736 N$21472 N$21471 "Straight Waveguide" sch_x=-223 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10737 N$21474 N$21473 "Straight Waveguide" sch_x=-221 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10738 N$21476 N$21475 "Straight Waveguide" sch_x=-221 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10739 N$21478 N$21477 "Straight Waveguide" sch_x=-221 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10740 N$21480 N$21479 "Straight Waveguide" sch_x=-221 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10741 N$21482 N$21481 "Straight Waveguide" sch_x=-221 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10742 N$21484 N$21483 "Straight Waveguide" sch_x=-221 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10743 N$21486 N$21485 "Straight Waveguide" sch_x=-221 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10744 N$21488 N$21487 "Straight Waveguide" sch_x=-221 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10745 N$21490 N$21489 "Straight Waveguide" sch_x=-221 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10746 N$21492 N$21491 "Straight Waveguide" sch_x=-221 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10747 N$21494 N$21493 "Straight Waveguide" sch_x=-221 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10748 N$21496 N$21495 "Straight Waveguide" sch_x=-221 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10749 N$21498 N$21497 "Straight Waveguide" sch_x=-221 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10750 N$21500 N$21499 "Straight Waveguide" sch_x=-221 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10751 N$21502 N$21501 "Straight Waveguide" sch_x=-221 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10752 N$21504 N$21503 "Straight Waveguide" sch_x=-221 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10753 N$21506 N$21505 "Straight Waveguide" sch_x=-221 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10754 N$21508 N$21507 "Straight Waveguide" sch_x=-221 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10755 N$21510 N$21509 "Straight Waveguide" sch_x=-221 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10756 N$21512 N$21511 "Straight Waveguide" sch_x=-221 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10757 N$21514 N$21513 "Straight Waveguide" sch_x=-221 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10758 N$21516 N$21515 "Straight Waveguide" sch_x=-221 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10759 N$21518 N$21517 "Straight Waveguide" sch_x=-221 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10760 N$21520 N$21519 "Straight Waveguide" sch_x=-221 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10761 N$21522 N$21521 "Straight Waveguide" sch_x=-221 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10762 N$21524 N$21523 "Straight Waveguide" sch_x=-221 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10763 N$21526 N$21525 "Straight Waveguide" sch_x=-221 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10764 N$21528 N$21527 "Straight Waveguide" sch_x=-221 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10765 N$21530 N$21529 "Straight Waveguide" sch_x=-221 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10766 N$21532 N$21531 "Straight Waveguide" sch_x=-221 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10767 N$21534 N$21533 "Straight Waveguide" sch_x=-221 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10768 N$21536 N$21535 "Straight Waveguide" sch_x=-221 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10769 N$21538 N$21537 "Straight Waveguide" sch_x=-221 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10770 N$21540 N$21539 "Straight Waveguide" sch_x=-221 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10771 N$21542 N$21541 "Straight Waveguide" sch_x=-221 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10772 N$21544 N$21543 "Straight Waveguide" sch_x=-221 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10773 N$21546 N$21545 "Straight Waveguide" sch_x=-221 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10774 N$21548 N$21547 "Straight Waveguide" sch_x=-221 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10775 N$21550 N$21549 "Straight Waveguide" sch_x=-221 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10776 N$21552 N$21551 "Straight Waveguide" sch_x=-221 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10777 N$21554 N$21553 "Straight Waveguide" sch_x=-221 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10778 N$21556 N$21555 "Straight Waveguide" sch_x=-221 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10779 N$21558 N$21557 "Straight Waveguide" sch_x=-221 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10780 N$21560 N$21559 "Straight Waveguide" sch_x=-221 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10781 N$21562 N$21561 "Straight Waveguide" sch_x=-221 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10782 N$21564 N$21563 "Straight Waveguide" sch_x=-221 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10783 N$21566 N$21565 "Straight Waveguide" sch_x=-221 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10784 N$21568 N$21567 "Straight Waveguide" sch_x=-221 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10785 N$21570 N$21569 "Straight Waveguide" sch_x=-221 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10786 N$21572 N$21571 "Straight Waveguide" sch_x=-221 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10787 N$21574 N$21573 "Straight Waveguide" sch_x=-221 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10788 N$21576 N$21575 "Straight Waveguide" sch_x=-221 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10789 N$21578 N$21577 "Straight Waveguide" sch_x=-221 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10790 N$21580 N$21579 "Straight Waveguide" sch_x=-221 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10791 N$21582 N$21581 "Straight Waveguide" sch_x=-221 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10792 N$21584 N$21583 "Straight Waveguide" sch_x=-221 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10793 N$21586 N$21585 "Straight Waveguide" sch_x=-221 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10794 N$21588 N$21587 "Straight Waveguide" sch_x=-221 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10795 N$21590 N$21589 "Straight Waveguide" sch_x=-221 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10796 N$21592 N$21591 "Straight Waveguide" sch_x=-221 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10797 N$21594 N$21593 "Straight Waveguide" sch_x=-221 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10798 N$21596 N$21595 "Straight Waveguide" sch_x=-221 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10799 N$21598 N$21597 "Straight Waveguide" sch_x=-221 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10800 N$21600 N$21599 "Straight Waveguide" sch_x=-221 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10801 N$21602 N$21601 "Straight Waveguide" sch_x=-221 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10802 N$21604 N$21603 "Straight Waveguide" sch_x=-221 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10803 N$21606 N$21605 "Straight Waveguide" sch_x=-221 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10804 N$21608 N$21607 "Straight Waveguide" sch_x=-221 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10805 N$21610 N$21609 "Straight Waveguide" sch_x=-221 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10806 N$21612 N$21611 "Straight Waveguide" sch_x=-221 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10807 N$21614 N$21613 "Straight Waveguide" sch_x=-221 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10808 N$21616 N$21615 "Straight Waveguide" sch_x=-221 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10809 N$21618 N$21617 "Straight Waveguide" sch_x=-221 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10810 N$21620 N$21619 "Straight Waveguide" sch_x=-221 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10811 N$21622 N$21621 "Straight Waveguide" sch_x=-221 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10812 N$21624 N$21623 "Straight Waveguide" sch_x=-221 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10813 N$21626 N$21625 "Straight Waveguide" sch_x=-221 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10814 N$21628 N$21627 "Straight Waveguide" sch_x=-221 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10815 N$21630 N$21629 "Straight Waveguide" sch_x=-221 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10816 N$21632 N$21631 "Straight Waveguide" sch_x=-221 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10817 N$21634 N$21633 "Straight Waveguide" sch_x=-221 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10818 N$21636 N$21635 "Straight Waveguide" sch_x=-221 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10819 N$21638 N$21637 "Straight Waveguide" sch_x=-221 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10820 N$21640 N$21639 "Straight Waveguide" sch_x=-221 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10821 N$21642 N$21641 "Straight Waveguide" sch_x=-221 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10822 N$21644 N$21643 "Straight Waveguide" sch_x=-221 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10823 N$21646 N$21645 "Straight Waveguide" sch_x=-221 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10824 N$21648 N$21647 "Straight Waveguide" sch_x=-221 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10825 N$21650 N$21649 "Straight Waveguide" sch_x=-221 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10826 N$21652 N$21651 "Straight Waveguide" sch_x=-221 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10827 N$21654 N$21653 "Straight Waveguide" sch_x=-221 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10828 N$21656 N$21655 "Straight Waveguide" sch_x=-221 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10829 N$21658 N$21657 "Straight Waveguide" sch_x=-221 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10830 N$21660 N$21659 "Straight Waveguide" sch_x=-221 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10831 N$21662 N$21661 "Straight Waveguide" sch_x=-219 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10832 N$21664 N$21663 "Straight Waveguide" sch_x=-219 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10833 N$21666 N$21665 "Straight Waveguide" sch_x=-219 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10834 N$21668 N$21667 "Straight Waveguide" sch_x=-219 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10835 N$21670 N$21669 "Straight Waveguide" sch_x=-219 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10836 N$21672 N$21671 "Straight Waveguide" sch_x=-219 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10837 N$21674 N$21673 "Straight Waveguide" sch_x=-219 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10838 N$21676 N$21675 "Straight Waveguide" sch_x=-219 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10839 N$21678 N$21677 "Straight Waveguide" sch_x=-219 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10840 N$21680 N$21679 "Straight Waveguide" sch_x=-219 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10841 N$21682 N$21681 "Straight Waveguide" sch_x=-219 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10842 N$21684 N$21683 "Straight Waveguide" sch_x=-219 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10843 N$21686 N$21685 "Straight Waveguide" sch_x=-219 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10844 N$21688 N$21687 "Straight Waveguide" sch_x=-219 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10845 N$21690 N$21689 "Straight Waveguide" sch_x=-219 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10846 N$21692 N$21691 "Straight Waveguide" sch_x=-219 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10847 N$21694 N$21693 "Straight Waveguide" sch_x=-219 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10848 N$21696 N$21695 "Straight Waveguide" sch_x=-219 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10849 N$21698 N$21697 "Straight Waveguide" sch_x=-219 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10850 N$21700 N$21699 "Straight Waveguide" sch_x=-219 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10851 N$21702 N$21701 "Straight Waveguide" sch_x=-219 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10852 N$21704 N$21703 "Straight Waveguide" sch_x=-219 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10853 N$21706 N$21705 "Straight Waveguide" sch_x=-219 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10854 N$21708 N$21707 "Straight Waveguide" sch_x=-219 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10855 N$21710 N$21709 "Straight Waveguide" sch_x=-219 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10856 N$21712 N$21711 "Straight Waveguide" sch_x=-219 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10857 N$21714 N$21713 "Straight Waveguide" sch_x=-219 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10858 N$21716 N$21715 "Straight Waveguide" sch_x=-219 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10859 N$21718 N$21717 "Straight Waveguide" sch_x=-219 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10860 N$21720 N$21719 "Straight Waveguide" sch_x=-219 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10861 N$21722 N$21721 "Straight Waveguide" sch_x=-219 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10862 N$21724 N$21723 "Straight Waveguide" sch_x=-219 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10863 N$21726 N$21725 "Straight Waveguide" sch_x=-219 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10864 N$21728 N$21727 "Straight Waveguide" sch_x=-219 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10865 N$21730 N$21729 "Straight Waveguide" sch_x=-219 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10866 N$21732 N$21731 "Straight Waveguide" sch_x=-219 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10867 N$21734 N$21733 "Straight Waveguide" sch_x=-219 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10868 N$21736 N$21735 "Straight Waveguide" sch_x=-219 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10869 N$21738 N$21737 "Straight Waveguide" sch_x=-219 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10870 N$21740 N$21739 "Straight Waveguide" sch_x=-219 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10871 N$21742 N$21741 "Straight Waveguide" sch_x=-219 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10872 N$21744 N$21743 "Straight Waveguide" sch_x=-219 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10873 N$21746 N$21745 "Straight Waveguide" sch_x=-219 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10874 N$21748 N$21747 "Straight Waveguide" sch_x=-219 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10875 N$21750 N$21749 "Straight Waveguide" sch_x=-219 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10876 N$21752 N$21751 "Straight Waveguide" sch_x=-219 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10877 N$21754 N$21753 "Straight Waveguide" sch_x=-219 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10878 N$21756 N$21755 "Straight Waveguide" sch_x=-219 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10879 N$21758 N$21757 "Straight Waveguide" sch_x=-219 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10880 N$21760 N$21759 "Straight Waveguide" sch_x=-219 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10881 N$21762 N$21761 "Straight Waveguide" sch_x=-219 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10882 N$21764 N$21763 "Straight Waveguide" sch_x=-219 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10883 N$21766 N$21765 "Straight Waveguide" sch_x=-219 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10884 N$21768 N$21767 "Straight Waveguide" sch_x=-219 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10885 N$21770 N$21769 "Straight Waveguide" sch_x=-219 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10886 N$21772 N$21771 "Straight Waveguide" sch_x=-219 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10887 N$21774 N$21773 "Straight Waveguide" sch_x=-219 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10888 N$21776 N$21775 "Straight Waveguide" sch_x=-219 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10889 N$21778 N$21777 "Straight Waveguide" sch_x=-219 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10890 N$21780 N$21779 "Straight Waveguide" sch_x=-219 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10891 N$21782 N$21781 "Straight Waveguide" sch_x=-219 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10892 N$21784 N$21783 "Straight Waveguide" sch_x=-219 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10893 N$21786 N$21785 "Straight Waveguide" sch_x=-219 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10894 N$21788 N$21787 "Straight Waveguide" sch_x=-219 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10895 N$21790 N$21789 "Straight Waveguide" sch_x=-219 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10896 N$21792 N$21791 "Straight Waveguide" sch_x=-219 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10897 N$21794 N$21793 "Straight Waveguide" sch_x=-219 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10898 N$21796 N$21795 "Straight Waveguide" sch_x=-219 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10899 N$21798 N$21797 "Straight Waveguide" sch_x=-219 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10900 N$21800 N$21799 "Straight Waveguide" sch_x=-219 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10901 N$21802 N$21801 "Straight Waveguide" sch_x=-219 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10902 N$21804 N$21803 "Straight Waveguide" sch_x=-219 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10903 N$21806 N$21805 "Straight Waveguide" sch_x=-219 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10904 N$21808 N$21807 "Straight Waveguide" sch_x=-219 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10905 N$21810 N$21809 "Straight Waveguide" sch_x=-219 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10906 N$21812 N$21811 "Straight Waveguide" sch_x=-219 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10907 N$21814 N$21813 "Straight Waveguide" sch_x=-219 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10908 N$21816 N$21815 "Straight Waveguide" sch_x=-219 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10909 N$21818 N$21817 "Straight Waveguide" sch_x=-219 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10910 N$21820 N$21819 "Straight Waveguide" sch_x=-219 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10911 N$21822 N$21821 "Straight Waveguide" sch_x=-219 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10912 N$21824 N$21823 "Straight Waveguide" sch_x=-219 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10913 N$21826 N$21825 "Straight Waveguide" sch_x=-219 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10914 N$21828 N$21827 "Straight Waveguide" sch_x=-219 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10915 N$21830 N$21829 "Straight Waveguide" sch_x=-219 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10916 N$21832 N$21831 "Straight Waveguide" sch_x=-219 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10917 N$21834 N$21833 "Straight Waveguide" sch_x=-219 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10918 N$21836 N$21835 "Straight Waveguide" sch_x=-219 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10919 N$21838 N$21837 "Straight Waveguide" sch_x=-219 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10920 N$21840 N$21839 "Straight Waveguide" sch_x=-219 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10921 N$21842 N$21841 "Straight Waveguide" sch_x=-219 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10922 N$21844 N$21843 "Straight Waveguide" sch_x=-219 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10923 N$21846 N$21845 "Straight Waveguide" sch_x=-217 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10924 N$21848 N$21847 "Straight Waveguide" sch_x=-217 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10925 N$21850 N$21849 "Straight Waveguide" sch_x=-217 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10926 N$21852 N$21851 "Straight Waveguide" sch_x=-217 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10927 N$21854 N$21853 "Straight Waveguide" sch_x=-217 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10928 N$21856 N$21855 "Straight Waveguide" sch_x=-217 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10929 N$21858 N$21857 "Straight Waveguide" sch_x=-217 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10930 N$21860 N$21859 "Straight Waveguide" sch_x=-217 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10931 N$21862 N$21861 "Straight Waveguide" sch_x=-217 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10932 N$21864 N$21863 "Straight Waveguide" sch_x=-217 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10933 N$21866 N$21865 "Straight Waveguide" sch_x=-217 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10934 N$21868 N$21867 "Straight Waveguide" sch_x=-217 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10935 N$21870 N$21869 "Straight Waveguide" sch_x=-217 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10936 N$21872 N$21871 "Straight Waveguide" sch_x=-217 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10937 N$21874 N$21873 "Straight Waveguide" sch_x=-217 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10938 N$21876 N$21875 "Straight Waveguide" sch_x=-217 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10939 N$21878 N$21877 "Straight Waveguide" sch_x=-217 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10940 N$21880 N$21879 "Straight Waveguide" sch_x=-217 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10941 N$21882 N$21881 "Straight Waveguide" sch_x=-217 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10942 N$21884 N$21883 "Straight Waveguide" sch_x=-217 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10943 N$21886 N$21885 "Straight Waveguide" sch_x=-217 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10944 N$21888 N$21887 "Straight Waveguide" sch_x=-217 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10945 N$21890 N$21889 "Straight Waveguide" sch_x=-217 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10946 N$21892 N$21891 "Straight Waveguide" sch_x=-217 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10947 N$21894 N$21893 "Straight Waveguide" sch_x=-217 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10948 N$21896 N$21895 "Straight Waveguide" sch_x=-217 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10949 N$21898 N$21897 "Straight Waveguide" sch_x=-217 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10950 N$21900 N$21899 "Straight Waveguide" sch_x=-217 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10951 N$21902 N$21901 "Straight Waveguide" sch_x=-217 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10952 N$21904 N$21903 "Straight Waveguide" sch_x=-217 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10953 N$21906 N$21905 "Straight Waveguide" sch_x=-217 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10954 N$21908 N$21907 "Straight Waveguide" sch_x=-217 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10955 N$21910 N$21909 "Straight Waveguide" sch_x=-217 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10956 N$21912 N$21911 "Straight Waveguide" sch_x=-217 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10957 N$21914 N$21913 "Straight Waveguide" sch_x=-217 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10958 N$21916 N$21915 "Straight Waveguide" sch_x=-217 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10959 N$21918 N$21917 "Straight Waveguide" sch_x=-217 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10960 N$21920 N$21919 "Straight Waveguide" sch_x=-217 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10961 N$21922 N$21921 "Straight Waveguide" sch_x=-217 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10962 N$21924 N$21923 "Straight Waveguide" sch_x=-217 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10963 N$21926 N$21925 "Straight Waveguide" sch_x=-217 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10964 N$21928 N$21927 "Straight Waveguide" sch_x=-217 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10965 N$21930 N$21929 "Straight Waveguide" sch_x=-217 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10966 N$21932 N$21931 "Straight Waveguide" sch_x=-217 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10967 N$21934 N$21933 "Straight Waveguide" sch_x=-217 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10968 N$21936 N$21935 "Straight Waveguide" sch_x=-217 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10969 N$21938 N$21937 "Straight Waveguide" sch_x=-217 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10970 N$21940 N$21939 "Straight Waveguide" sch_x=-217 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10971 N$21942 N$21941 "Straight Waveguide" sch_x=-217 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10972 N$21944 N$21943 "Straight Waveguide" sch_x=-217 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10973 N$21946 N$21945 "Straight Waveguide" sch_x=-217 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10974 N$21948 N$21947 "Straight Waveguide" sch_x=-217 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10975 N$21950 N$21949 "Straight Waveguide" sch_x=-217 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10976 N$21952 N$21951 "Straight Waveguide" sch_x=-217 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10977 N$21954 N$21953 "Straight Waveguide" sch_x=-217 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10978 N$21956 N$21955 "Straight Waveguide" sch_x=-217 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10979 N$21958 N$21957 "Straight Waveguide" sch_x=-217 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10980 N$21960 N$21959 "Straight Waveguide" sch_x=-217 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10981 N$21962 N$21961 "Straight Waveguide" sch_x=-217 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10982 N$21964 N$21963 "Straight Waveguide" sch_x=-217 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10983 N$21966 N$21965 "Straight Waveguide" sch_x=-217 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10984 N$21968 N$21967 "Straight Waveguide" sch_x=-217 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10985 N$21970 N$21969 "Straight Waveguide" sch_x=-217 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10986 N$21972 N$21971 "Straight Waveguide" sch_x=-217 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10987 N$21974 N$21973 "Straight Waveguide" sch_x=-217 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10988 N$21976 N$21975 "Straight Waveguide" sch_x=-217 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10989 N$21978 N$21977 "Straight Waveguide" sch_x=-217 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10990 N$21980 N$21979 "Straight Waveguide" sch_x=-217 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10991 N$21982 N$21981 "Straight Waveguide" sch_x=-217 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10992 N$21984 N$21983 "Straight Waveguide" sch_x=-217 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10993 N$21986 N$21985 "Straight Waveguide" sch_x=-217 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10994 N$21988 N$21987 "Straight Waveguide" sch_x=-217 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10995 N$21990 N$21989 "Straight Waveguide" sch_x=-217 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10996 N$21992 N$21991 "Straight Waveguide" sch_x=-217 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10997 N$21994 N$21993 "Straight Waveguide" sch_x=-217 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10998 N$21996 N$21995 "Straight Waveguide" sch_x=-217 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10999 N$21998 N$21997 "Straight Waveguide" sch_x=-217 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11000 N$22000 N$21999 "Straight Waveguide" sch_x=-217 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11001 N$22002 N$22001 "Straight Waveguide" sch_x=-217 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11002 N$22004 N$22003 "Straight Waveguide" sch_x=-217 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11003 N$22006 N$22005 "Straight Waveguide" sch_x=-217 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11004 N$22008 N$22007 "Straight Waveguide" sch_x=-217 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11005 N$22010 N$22009 "Straight Waveguide" sch_x=-217 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11006 N$22012 N$22011 "Straight Waveguide" sch_x=-217 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11007 N$22014 N$22013 "Straight Waveguide" sch_x=-217 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11008 N$22016 N$22015 "Straight Waveguide" sch_x=-217 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11009 N$22018 N$22017 "Straight Waveguide" sch_x=-217 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11010 N$22020 N$22019 "Straight Waveguide" sch_x=-217 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11011 N$22022 N$22021 "Straight Waveguide" sch_x=-217 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11012 N$22024 N$22023 "Straight Waveguide" sch_x=-217 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11013 N$22026 N$22025 "Straight Waveguide" sch_x=-215 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11014 N$22028 N$22027 "Straight Waveguide" sch_x=-215 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11015 N$22030 N$22029 "Straight Waveguide" sch_x=-215 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11016 N$22032 N$22031 "Straight Waveguide" sch_x=-215 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11017 N$22034 N$22033 "Straight Waveguide" sch_x=-215 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11018 N$22036 N$22035 "Straight Waveguide" sch_x=-215 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11019 N$22038 N$22037 "Straight Waveguide" sch_x=-215 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11020 N$22040 N$22039 "Straight Waveguide" sch_x=-215 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11021 N$22042 N$22041 "Straight Waveguide" sch_x=-215 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11022 N$22044 N$22043 "Straight Waveguide" sch_x=-215 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11023 N$22046 N$22045 "Straight Waveguide" sch_x=-215 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11024 N$22048 N$22047 "Straight Waveguide" sch_x=-215 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11025 N$22050 N$22049 "Straight Waveguide" sch_x=-215 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11026 N$22052 N$22051 "Straight Waveguide" sch_x=-215 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11027 N$22054 N$22053 "Straight Waveguide" sch_x=-215 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11028 N$22056 N$22055 "Straight Waveguide" sch_x=-215 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11029 N$22058 N$22057 "Straight Waveguide" sch_x=-215 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11030 N$22060 N$22059 "Straight Waveguide" sch_x=-215 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11031 N$22062 N$22061 "Straight Waveguide" sch_x=-215 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11032 N$22064 N$22063 "Straight Waveguide" sch_x=-215 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11033 N$22066 N$22065 "Straight Waveguide" sch_x=-215 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11034 N$22068 N$22067 "Straight Waveguide" sch_x=-215 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11035 N$22070 N$22069 "Straight Waveguide" sch_x=-215 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11036 N$22072 N$22071 "Straight Waveguide" sch_x=-215 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11037 N$22074 N$22073 "Straight Waveguide" sch_x=-215 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11038 N$22076 N$22075 "Straight Waveguide" sch_x=-215 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11039 N$22078 N$22077 "Straight Waveguide" sch_x=-215 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11040 N$22080 N$22079 "Straight Waveguide" sch_x=-215 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11041 N$22082 N$22081 "Straight Waveguide" sch_x=-215 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11042 N$22084 N$22083 "Straight Waveguide" sch_x=-215 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11043 N$22086 N$22085 "Straight Waveguide" sch_x=-215 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11044 N$22088 N$22087 "Straight Waveguide" sch_x=-215 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11045 N$22090 N$22089 "Straight Waveguide" sch_x=-215 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11046 N$22092 N$22091 "Straight Waveguide" sch_x=-215 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11047 N$22094 N$22093 "Straight Waveguide" sch_x=-215 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11048 N$22096 N$22095 "Straight Waveguide" sch_x=-215 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11049 N$22098 N$22097 "Straight Waveguide" sch_x=-215 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11050 N$22100 N$22099 "Straight Waveguide" sch_x=-215 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11051 N$22102 N$22101 "Straight Waveguide" sch_x=-215 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11052 N$22104 N$22103 "Straight Waveguide" sch_x=-215 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11053 N$22106 N$22105 "Straight Waveguide" sch_x=-215 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11054 N$22108 N$22107 "Straight Waveguide" sch_x=-215 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11055 N$22110 N$22109 "Straight Waveguide" sch_x=-215 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11056 N$22112 N$22111 "Straight Waveguide" sch_x=-215 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11057 N$22114 N$22113 "Straight Waveguide" sch_x=-215 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11058 N$22116 N$22115 "Straight Waveguide" sch_x=-215 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11059 N$22118 N$22117 "Straight Waveguide" sch_x=-215 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11060 N$22120 N$22119 "Straight Waveguide" sch_x=-215 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11061 N$22122 N$22121 "Straight Waveguide" sch_x=-215 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11062 N$22124 N$22123 "Straight Waveguide" sch_x=-215 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11063 N$22126 N$22125 "Straight Waveguide" sch_x=-215 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11064 N$22128 N$22127 "Straight Waveguide" sch_x=-215 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11065 N$22130 N$22129 "Straight Waveguide" sch_x=-215 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11066 N$22132 N$22131 "Straight Waveguide" sch_x=-215 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11067 N$22134 N$22133 "Straight Waveguide" sch_x=-215 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11068 N$22136 N$22135 "Straight Waveguide" sch_x=-215 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11069 N$22138 N$22137 "Straight Waveguide" sch_x=-215 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11070 N$22140 N$22139 "Straight Waveguide" sch_x=-215 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11071 N$22142 N$22141 "Straight Waveguide" sch_x=-215 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11072 N$22144 N$22143 "Straight Waveguide" sch_x=-215 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11073 N$22146 N$22145 "Straight Waveguide" sch_x=-215 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11074 N$22148 N$22147 "Straight Waveguide" sch_x=-215 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11075 N$22150 N$22149 "Straight Waveguide" sch_x=-215 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11076 N$22152 N$22151 "Straight Waveguide" sch_x=-215 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11077 N$22154 N$22153 "Straight Waveguide" sch_x=-215 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11078 N$22156 N$22155 "Straight Waveguide" sch_x=-215 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11079 N$22158 N$22157 "Straight Waveguide" sch_x=-215 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11080 N$22160 N$22159 "Straight Waveguide" sch_x=-215 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11081 N$22162 N$22161 "Straight Waveguide" sch_x=-215 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11082 N$22164 N$22163 "Straight Waveguide" sch_x=-215 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11083 N$22166 N$22165 "Straight Waveguide" sch_x=-215 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11084 N$22168 N$22167 "Straight Waveguide" sch_x=-215 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11085 N$22170 N$22169 "Straight Waveguide" sch_x=-215 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11086 N$22172 N$22171 "Straight Waveguide" sch_x=-215 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11087 N$22174 N$22173 "Straight Waveguide" sch_x=-215 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11088 N$22176 N$22175 "Straight Waveguide" sch_x=-215 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11089 N$22178 N$22177 "Straight Waveguide" sch_x=-215 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11090 N$22180 N$22179 "Straight Waveguide" sch_x=-215 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11091 N$22182 N$22181 "Straight Waveguide" sch_x=-215 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11092 N$22184 N$22183 "Straight Waveguide" sch_x=-215 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11093 N$22186 N$22185 "Straight Waveguide" sch_x=-215 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11094 N$22188 N$22187 "Straight Waveguide" sch_x=-215 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11095 N$22190 N$22189 "Straight Waveguide" sch_x=-215 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11096 N$22192 N$22191 "Straight Waveguide" sch_x=-215 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11097 N$22194 N$22193 "Straight Waveguide" sch_x=-215 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11098 N$22196 N$22195 "Straight Waveguide" sch_x=-215 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11099 N$22198 N$22197 "Straight Waveguide" sch_x=-215 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11100 N$22200 N$22199 "Straight Waveguide" sch_x=-215 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11101 N$22202 N$22201 "Straight Waveguide" sch_x=-213 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11102 N$22204 N$22203 "Straight Waveguide" sch_x=-213 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11103 N$22206 N$22205 "Straight Waveguide" sch_x=-213 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11104 N$22208 N$22207 "Straight Waveguide" sch_x=-213 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11105 N$22210 N$22209 "Straight Waveguide" sch_x=-213 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11106 N$22212 N$22211 "Straight Waveguide" sch_x=-213 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11107 N$22214 N$22213 "Straight Waveguide" sch_x=-213 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11108 N$22216 N$22215 "Straight Waveguide" sch_x=-213 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11109 N$22218 N$22217 "Straight Waveguide" sch_x=-213 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11110 N$22220 N$22219 "Straight Waveguide" sch_x=-213 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11111 N$22222 N$22221 "Straight Waveguide" sch_x=-213 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11112 N$22224 N$22223 "Straight Waveguide" sch_x=-213 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11113 N$22226 N$22225 "Straight Waveguide" sch_x=-213 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11114 N$22228 N$22227 "Straight Waveguide" sch_x=-213 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11115 N$22230 N$22229 "Straight Waveguide" sch_x=-213 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11116 N$22232 N$22231 "Straight Waveguide" sch_x=-213 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11117 N$22234 N$22233 "Straight Waveguide" sch_x=-213 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11118 N$22236 N$22235 "Straight Waveguide" sch_x=-213 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11119 N$22238 N$22237 "Straight Waveguide" sch_x=-213 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11120 N$22240 N$22239 "Straight Waveguide" sch_x=-213 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11121 N$22242 N$22241 "Straight Waveguide" sch_x=-213 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11122 N$22244 N$22243 "Straight Waveguide" sch_x=-213 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11123 N$22246 N$22245 "Straight Waveguide" sch_x=-213 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11124 N$22248 N$22247 "Straight Waveguide" sch_x=-213 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11125 N$22250 N$22249 "Straight Waveguide" sch_x=-213 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11126 N$22252 N$22251 "Straight Waveguide" sch_x=-213 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11127 N$22254 N$22253 "Straight Waveguide" sch_x=-213 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11128 N$22256 N$22255 "Straight Waveguide" sch_x=-213 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11129 N$22258 N$22257 "Straight Waveguide" sch_x=-213 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11130 N$22260 N$22259 "Straight Waveguide" sch_x=-213 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11131 N$22262 N$22261 "Straight Waveguide" sch_x=-213 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11132 N$22264 N$22263 "Straight Waveguide" sch_x=-213 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11133 N$22266 N$22265 "Straight Waveguide" sch_x=-213 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11134 N$22268 N$22267 "Straight Waveguide" sch_x=-213 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11135 N$22270 N$22269 "Straight Waveguide" sch_x=-213 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11136 N$22272 N$22271 "Straight Waveguide" sch_x=-213 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11137 N$22274 N$22273 "Straight Waveguide" sch_x=-213 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11138 N$22276 N$22275 "Straight Waveguide" sch_x=-213 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11139 N$22278 N$22277 "Straight Waveguide" sch_x=-213 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11140 N$22280 N$22279 "Straight Waveguide" sch_x=-213 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11141 N$22282 N$22281 "Straight Waveguide" sch_x=-213 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11142 N$22284 N$22283 "Straight Waveguide" sch_x=-213 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11143 N$22286 N$22285 "Straight Waveguide" sch_x=-213 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11144 N$22288 N$22287 "Straight Waveguide" sch_x=-213 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11145 N$22290 N$22289 "Straight Waveguide" sch_x=-213 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11146 N$22292 N$22291 "Straight Waveguide" sch_x=-213 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11147 N$22294 N$22293 "Straight Waveguide" sch_x=-213 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11148 N$22296 N$22295 "Straight Waveguide" sch_x=-213 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11149 N$22298 N$22297 "Straight Waveguide" sch_x=-213 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11150 N$22300 N$22299 "Straight Waveguide" sch_x=-213 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11151 N$22302 N$22301 "Straight Waveguide" sch_x=-213 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11152 N$22304 N$22303 "Straight Waveguide" sch_x=-213 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11153 N$22306 N$22305 "Straight Waveguide" sch_x=-213 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11154 N$22308 N$22307 "Straight Waveguide" sch_x=-213 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11155 N$22310 N$22309 "Straight Waveguide" sch_x=-213 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11156 N$22312 N$22311 "Straight Waveguide" sch_x=-213 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11157 N$22314 N$22313 "Straight Waveguide" sch_x=-213 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11158 N$22316 N$22315 "Straight Waveguide" sch_x=-213 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11159 N$22318 N$22317 "Straight Waveguide" sch_x=-213 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11160 N$22320 N$22319 "Straight Waveguide" sch_x=-213 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11161 N$22322 N$22321 "Straight Waveguide" sch_x=-213 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11162 N$22324 N$22323 "Straight Waveguide" sch_x=-213 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11163 N$22326 N$22325 "Straight Waveguide" sch_x=-213 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11164 N$22328 N$22327 "Straight Waveguide" sch_x=-213 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11165 N$22330 N$22329 "Straight Waveguide" sch_x=-213 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11166 N$22332 N$22331 "Straight Waveguide" sch_x=-213 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11167 N$22334 N$22333 "Straight Waveguide" sch_x=-213 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11168 N$22336 N$22335 "Straight Waveguide" sch_x=-213 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11169 N$22338 N$22337 "Straight Waveguide" sch_x=-213 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11170 N$22340 N$22339 "Straight Waveguide" sch_x=-213 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11171 N$22342 N$22341 "Straight Waveguide" sch_x=-213 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11172 N$22344 N$22343 "Straight Waveguide" sch_x=-213 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11173 N$22346 N$22345 "Straight Waveguide" sch_x=-213 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11174 N$22348 N$22347 "Straight Waveguide" sch_x=-213 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11175 N$22350 N$22349 "Straight Waveguide" sch_x=-213 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11176 N$22352 N$22351 "Straight Waveguide" sch_x=-213 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11177 N$22354 N$22353 "Straight Waveguide" sch_x=-213 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11178 N$22356 N$22355 "Straight Waveguide" sch_x=-213 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11179 N$22358 N$22357 "Straight Waveguide" sch_x=-213 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11180 N$22360 N$22359 "Straight Waveguide" sch_x=-213 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11181 N$22362 N$22361 "Straight Waveguide" sch_x=-213 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11182 N$22364 N$22363 "Straight Waveguide" sch_x=-213 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11183 N$22366 N$22365 "Straight Waveguide" sch_x=-213 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11184 N$22368 N$22367 "Straight Waveguide" sch_x=-213 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11185 N$22370 N$22369 "Straight Waveguide" sch_x=-213 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11186 N$22372 N$22371 "Straight Waveguide" sch_x=-213 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11187 N$22374 N$22373 "Straight Waveguide" sch_x=-211 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11188 N$22376 N$22375 "Straight Waveguide" sch_x=-211 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11189 N$22378 N$22377 "Straight Waveguide" sch_x=-211 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11190 N$22380 N$22379 "Straight Waveguide" sch_x=-211 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11191 N$22382 N$22381 "Straight Waveguide" sch_x=-211 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11192 N$22384 N$22383 "Straight Waveguide" sch_x=-211 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11193 N$22386 N$22385 "Straight Waveguide" sch_x=-211 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11194 N$22388 N$22387 "Straight Waveguide" sch_x=-211 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11195 N$22390 N$22389 "Straight Waveguide" sch_x=-211 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11196 N$22392 N$22391 "Straight Waveguide" sch_x=-211 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11197 N$22394 N$22393 "Straight Waveguide" sch_x=-211 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11198 N$22396 N$22395 "Straight Waveguide" sch_x=-211 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11199 N$22398 N$22397 "Straight Waveguide" sch_x=-211 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11200 N$22400 N$22399 "Straight Waveguide" sch_x=-211 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11201 N$22402 N$22401 "Straight Waveguide" sch_x=-211 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11202 N$22404 N$22403 "Straight Waveguide" sch_x=-211 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11203 N$22406 N$22405 "Straight Waveguide" sch_x=-211 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11204 N$22408 N$22407 "Straight Waveguide" sch_x=-211 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11205 N$22410 N$22409 "Straight Waveguide" sch_x=-211 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11206 N$22412 N$22411 "Straight Waveguide" sch_x=-211 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11207 N$22414 N$22413 "Straight Waveguide" sch_x=-211 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11208 N$22416 N$22415 "Straight Waveguide" sch_x=-211 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11209 N$22418 N$22417 "Straight Waveguide" sch_x=-211 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11210 N$22420 N$22419 "Straight Waveguide" sch_x=-211 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11211 N$22422 N$22421 "Straight Waveguide" sch_x=-211 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11212 N$22424 N$22423 "Straight Waveguide" sch_x=-211 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11213 N$22426 N$22425 "Straight Waveguide" sch_x=-211 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11214 N$22428 N$22427 "Straight Waveguide" sch_x=-211 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11215 N$22430 N$22429 "Straight Waveguide" sch_x=-211 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11216 N$22432 N$22431 "Straight Waveguide" sch_x=-211 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11217 N$22434 N$22433 "Straight Waveguide" sch_x=-211 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11218 N$22436 N$22435 "Straight Waveguide" sch_x=-211 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11219 N$22438 N$22437 "Straight Waveguide" sch_x=-211 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11220 N$22440 N$22439 "Straight Waveguide" sch_x=-211 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11221 N$22442 N$22441 "Straight Waveguide" sch_x=-211 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11222 N$22444 N$22443 "Straight Waveguide" sch_x=-211 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11223 N$22446 N$22445 "Straight Waveguide" sch_x=-211 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11224 N$22448 N$22447 "Straight Waveguide" sch_x=-211 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11225 N$22450 N$22449 "Straight Waveguide" sch_x=-211 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11226 N$22452 N$22451 "Straight Waveguide" sch_x=-211 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11227 N$22454 N$22453 "Straight Waveguide" sch_x=-211 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11228 N$22456 N$22455 "Straight Waveguide" sch_x=-211 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11229 N$22458 N$22457 "Straight Waveguide" sch_x=-211 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11230 N$22460 N$22459 "Straight Waveguide" sch_x=-211 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11231 N$22462 N$22461 "Straight Waveguide" sch_x=-211 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11232 N$22464 N$22463 "Straight Waveguide" sch_x=-211 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11233 N$22466 N$22465 "Straight Waveguide" sch_x=-211 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11234 N$22468 N$22467 "Straight Waveguide" sch_x=-211 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11235 N$22470 N$22469 "Straight Waveguide" sch_x=-211 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11236 N$22472 N$22471 "Straight Waveguide" sch_x=-211 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11237 N$22474 N$22473 "Straight Waveguide" sch_x=-211 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11238 N$22476 N$22475 "Straight Waveguide" sch_x=-211 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11239 N$22478 N$22477 "Straight Waveguide" sch_x=-211 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11240 N$22480 N$22479 "Straight Waveguide" sch_x=-211 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11241 N$22482 N$22481 "Straight Waveguide" sch_x=-211 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11242 N$22484 N$22483 "Straight Waveguide" sch_x=-211 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11243 N$22486 N$22485 "Straight Waveguide" sch_x=-211 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11244 N$22488 N$22487 "Straight Waveguide" sch_x=-211 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11245 N$22490 N$22489 "Straight Waveguide" sch_x=-211 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11246 N$22492 N$22491 "Straight Waveguide" sch_x=-211 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11247 N$22494 N$22493 "Straight Waveguide" sch_x=-211 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11248 N$22496 N$22495 "Straight Waveguide" sch_x=-211 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11249 N$22498 N$22497 "Straight Waveguide" sch_x=-211 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11250 N$22500 N$22499 "Straight Waveguide" sch_x=-211 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11251 N$22502 N$22501 "Straight Waveguide" sch_x=-211 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11252 N$22504 N$22503 "Straight Waveguide" sch_x=-211 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11253 N$22506 N$22505 "Straight Waveguide" sch_x=-211 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11254 N$22508 N$22507 "Straight Waveguide" sch_x=-211 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11255 N$22510 N$22509 "Straight Waveguide" sch_x=-211 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11256 N$22512 N$22511 "Straight Waveguide" sch_x=-211 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11257 N$22514 N$22513 "Straight Waveguide" sch_x=-211 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11258 N$22516 N$22515 "Straight Waveguide" sch_x=-211 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11259 N$22518 N$22517 "Straight Waveguide" sch_x=-211 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11260 N$22520 N$22519 "Straight Waveguide" sch_x=-211 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11261 N$22522 N$22521 "Straight Waveguide" sch_x=-211 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11262 N$22524 N$22523 "Straight Waveguide" sch_x=-211 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11263 N$22526 N$22525 "Straight Waveguide" sch_x=-211 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11264 N$22528 N$22527 "Straight Waveguide" sch_x=-211 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11265 N$22530 N$22529 "Straight Waveguide" sch_x=-211 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11266 N$22532 N$22531 "Straight Waveguide" sch_x=-211 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11267 N$22534 N$22533 "Straight Waveguide" sch_x=-211 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11268 N$22536 N$22535 "Straight Waveguide" sch_x=-211 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11269 N$22538 N$22537 "Straight Waveguide" sch_x=-211 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11270 N$22540 N$22539 "Straight Waveguide" sch_x=-211 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11271 N$22542 N$22541 "Straight Waveguide" sch_x=-209 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11272 N$22544 N$22543 "Straight Waveguide" sch_x=-209 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11273 N$22546 N$22545 "Straight Waveguide" sch_x=-209 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11274 N$22548 N$22547 "Straight Waveguide" sch_x=-209 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11275 N$22550 N$22549 "Straight Waveguide" sch_x=-209 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11276 N$22552 N$22551 "Straight Waveguide" sch_x=-209 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11277 N$22554 N$22553 "Straight Waveguide" sch_x=-209 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11278 N$22556 N$22555 "Straight Waveguide" sch_x=-209 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11279 N$22558 N$22557 "Straight Waveguide" sch_x=-209 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11280 N$22560 N$22559 "Straight Waveguide" sch_x=-209 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11281 N$22562 N$22561 "Straight Waveguide" sch_x=-209 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11282 N$22564 N$22563 "Straight Waveguide" sch_x=-209 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11283 N$22566 N$22565 "Straight Waveguide" sch_x=-209 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11284 N$22568 N$22567 "Straight Waveguide" sch_x=-209 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11285 N$22570 N$22569 "Straight Waveguide" sch_x=-209 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11286 N$22572 N$22571 "Straight Waveguide" sch_x=-209 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11287 N$22574 N$22573 "Straight Waveguide" sch_x=-209 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11288 N$22576 N$22575 "Straight Waveguide" sch_x=-209 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11289 N$22578 N$22577 "Straight Waveguide" sch_x=-209 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11290 N$22580 N$22579 "Straight Waveguide" sch_x=-209 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11291 N$22582 N$22581 "Straight Waveguide" sch_x=-209 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11292 N$22584 N$22583 "Straight Waveguide" sch_x=-209 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11293 N$22586 N$22585 "Straight Waveguide" sch_x=-209 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11294 N$22588 N$22587 "Straight Waveguide" sch_x=-209 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11295 N$22590 N$22589 "Straight Waveguide" sch_x=-209 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11296 N$22592 N$22591 "Straight Waveguide" sch_x=-209 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11297 N$22594 N$22593 "Straight Waveguide" sch_x=-209 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11298 N$22596 N$22595 "Straight Waveguide" sch_x=-209 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11299 N$22598 N$22597 "Straight Waveguide" sch_x=-209 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11300 N$22600 N$22599 "Straight Waveguide" sch_x=-209 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11301 N$22602 N$22601 "Straight Waveguide" sch_x=-209 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11302 N$22604 N$22603 "Straight Waveguide" sch_x=-209 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11303 N$22606 N$22605 "Straight Waveguide" sch_x=-209 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11304 N$22608 N$22607 "Straight Waveguide" sch_x=-209 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11305 N$22610 N$22609 "Straight Waveguide" sch_x=-209 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11306 N$22612 N$22611 "Straight Waveguide" sch_x=-209 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11307 N$22614 N$22613 "Straight Waveguide" sch_x=-209 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11308 N$22616 N$22615 "Straight Waveguide" sch_x=-209 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11309 N$22618 N$22617 "Straight Waveguide" sch_x=-209 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11310 N$22620 N$22619 "Straight Waveguide" sch_x=-209 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11311 N$22622 N$22621 "Straight Waveguide" sch_x=-209 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11312 N$22624 N$22623 "Straight Waveguide" sch_x=-209 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11313 N$22626 N$22625 "Straight Waveguide" sch_x=-209 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11314 N$22628 N$22627 "Straight Waveguide" sch_x=-209 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11315 N$22630 N$22629 "Straight Waveguide" sch_x=-209 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11316 N$22632 N$22631 "Straight Waveguide" sch_x=-209 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11317 N$22634 N$22633 "Straight Waveguide" sch_x=-209 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11318 N$22636 N$22635 "Straight Waveguide" sch_x=-209 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11319 N$22638 N$22637 "Straight Waveguide" sch_x=-209 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11320 N$22640 N$22639 "Straight Waveguide" sch_x=-209 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11321 N$22642 N$22641 "Straight Waveguide" sch_x=-209 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11322 N$22644 N$22643 "Straight Waveguide" sch_x=-209 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11323 N$22646 N$22645 "Straight Waveguide" sch_x=-209 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11324 N$22648 N$22647 "Straight Waveguide" sch_x=-209 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11325 N$22650 N$22649 "Straight Waveguide" sch_x=-209 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11326 N$22652 N$22651 "Straight Waveguide" sch_x=-209 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11327 N$22654 N$22653 "Straight Waveguide" sch_x=-209 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11328 N$22656 N$22655 "Straight Waveguide" sch_x=-209 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11329 N$22658 N$22657 "Straight Waveguide" sch_x=-209 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11330 N$22660 N$22659 "Straight Waveguide" sch_x=-209 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11331 N$22662 N$22661 "Straight Waveguide" sch_x=-209 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11332 N$22664 N$22663 "Straight Waveguide" sch_x=-209 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11333 N$22666 N$22665 "Straight Waveguide" sch_x=-209 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11334 N$22668 N$22667 "Straight Waveguide" sch_x=-209 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11335 N$22670 N$22669 "Straight Waveguide" sch_x=-209 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11336 N$22672 N$22671 "Straight Waveguide" sch_x=-209 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11337 N$22674 N$22673 "Straight Waveguide" sch_x=-209 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11338 N$22676 N$22675 "Straight Waveguide" sch_x=-209 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11339 N$22678 N$22677 "Straight Waveguide" sch_x=-209 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11340 N$22680 N$22679 "Straight Waveguide" sch_x=-209 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11341 N$22682 N$22681 "Straight Waveguide" sch_x=-209 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11342 N$22684 N$22683 "Straight Waveguide" sch_x=-209 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11343 N$22686 N$22685 "Straight Waveguide" sch_x=-209 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11344 N$22688 N$22687 "Straight Waveguide" sch_x=-209 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11345 N$22690 N$22689 "Straight Waveguide" sch_x=-209 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11346 N$22692 N$22691 "Straight Waveguide" sch_x=-209 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11347 N$22694 N$22693 "Straight Waveguide" sch_x=-209 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11348 N$22696 N$22695 "Straight Waveguide" sch_x=-209 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11349 N$22698 N$22697 "Straight Waveguide" sch_x=-209 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11350 N$22700 N$22699 "Straight Waveguide" sch_x=-209 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11351 N$22702 N$22701 "Straight Waveguide" sch_x=-209 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11352 N$22704 N$22703 "Straight Waveguide" sch_x=-209 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11353 N$22706 N$22705 "Straight Waveguide" sch_x=-207 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11354 N$22708 N$22707 "Straight Waveguide" sch_x=-207 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11355 N$22710 N$22709 "Straight Waveguide" sch_x=-207 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11356 N$22712 N$22711 "Straight Waveguide" sch_x=-207 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11357 N$22714 N$22713 "Straight Waveguide" sch_x=-207 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11358 N$22716 N$22715 "Straight Waveguide" sch_x=-207 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11359 N$22718 N$22717 "Straight Waveguide" sch_x=-207 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11360 N$22720 N$22719 "Straight Waveguide" sch_x=-207 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11361 N$22722 N$22721 "Straight Waveguide" sch_x=-207 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11362 N$22724 N$22723 "Straight Waveguide" sch_x=-207 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11363 N$22726 N$22725 "Straight Waveguide" sch_x=-207 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11364 N$22728 N$22727 "Straight Waveguide" sch_x=-207 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11365 N$22730 N$22729 "Straight Waveguide" sch_x=-207 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11366 N$22732 N$22731 "Straight Waveguide" sch_x=-207 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11367 N$22734 N$22733 "Straight Waveguide" sch_x=-207 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11368 N$22736 N$22735 "Straight Waveguide" sch_x=-207 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11369 N$22738 N$22737 "Straight Waveguide" sch_x=-207 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11370 N$22740 N$22739 "Straight Waveguide" sch_x=-207 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11371 N$22742 N$22741 "Straight Waveguide" sch_x=-207 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11372 N$22744 N$22743 "Straight Waveguide" sch_x=-207 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11373 N$22746 N$22745 "Straight Waveguide" sch_x=-207 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11374 N$22748 N$22747 "Straight Waveguide" sch_x=-207 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11375 N$22750 N$22749 "Straight Waveguide" sch_x=-207 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11376 N$22752 N$22751 "Straight Waveguide" sch_x=-207 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11377 N$22754 N$22753 "Straight Waveguide" sch_x=-207 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11378 N$22756 N$22755 "Straight Waveguide" sch_x=-207 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11379 N$22758 N$22757 "Straight Waveguide" sch_x=-207 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11380 N$22760 N$22759 "Straight Waveguide" sch_x=-207 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11381 N$22762 N$22761 "Straight Waveguide" sch_x=-207 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11382 N$22764 N$22763 "Straight Waveguide" sch_x=-207 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11383 N$22766 N$22765 "Straight Waveguide" sch_x=-207 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11384 N$22768 N$22767 "Straight Waveguide" sch_x=-207 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11385 N$22770 N$22769 "Straight Waveguide" sch_x=-207 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11386 N$22772 N$22771 "Straight Waveguide" sch_x=-207 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11387 N$22774 N$22773 "Straight Waveguide" sch_x=-207 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11388 N$22776 N$22775 "Straight Waveguide" sch_x=-207 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11389 N$22778 N$22777 "Straight Waveguide" sch_x=-207 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11390 N$22780 N$22779 "Straight Waveguide" sch_x=-207 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11391 N$22782 N$22781 "Straight Waveguide" sch_x=-207 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11392 N$22784 N$22783 "Straight Waveguide" sch_x=-207 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11393 N$22786 N$22785 "Straight Waveguide" sch_x=-207 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11394 N$22788 N$22787 "Straight Waveguide" sch_x=-207 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11395 N$22790 N$22789 "Straight Waveguide" sch_x=-207 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11396 N$22792 N$22791 "Straight Waveguide" sch_x=-207 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11397 N$22794 N$22793 "Straight Waveguide" sch_x=-207 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11398 N$22796 N$22795 "Straight Waveguide" sch_x=-207 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11399 N$22798 N$22797 "Straight Waveguide" sch_x=-207 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11400 N$22800 N$22799 "Straight Waveguide" sch_x=-207 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11401 N$22802 N$22801 "Straight Waveguide" sch_x=-207 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11402 N$22804 N$22803 "Straight Waveguide" sch_x=-207 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11403 N$22806 N$22805 "Straight Waveguide" sch_x=-207 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11404 N$22808 N$22807 "Straight Waveguide" sch_x=-207 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11405 N$22810 N$22809 "Straight Waveguide" sch_x=-207 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11406 N$22812 N$22811 "Straight Waveguide" sch_x=-207 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11407 N$22814 N$22813 "Straight Waveguide" sch_x=-207 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11408 N$22816 N$22815 "Straight Waveguide" sch_x=-207 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11409 N$22818 N$22817 "Straight Waveguide" sch_x=-207 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11410 N$22820 N$22819 "Straight Waveguide" sch_x=-207 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11411 N$22822 N$22821 "Straight Waveguide" sch_x=-207 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11412 N$22824 N$22823 "Straight Waveguide" sch_x=-207 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11413 N$22826 N$22825 "Straight Waveguide" sch_x=-207 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11414 N$22828 N$22827 "Straight Waveguide" sch_x=-207 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11415 N$22830 N$22829 "Straight Waveguide" sch_x=-207 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11416 N$22832 N$22831 "Straight Waveguide" sch_x=-207 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11417 N$22834 N$22833 "Straight Waveguide" sch_x=-207 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11418 N$22836 N$22835 "Straight Waveguide" sch_x=-207 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11419 N$22838 N$22837 "Straight Waveguide" sch_x=-207 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11420 N$22840 N$22839 "Straight Waveguide" sch_x=-207 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11421 N$22842 N$22841 "Straight Waveguide" sch_x=-207 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11422 N$22844 N$22843 "Straight Waveguide" sch_x=-207 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11423 N$22846 N$22845 "Straight Waveguide" sch_x=-207 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11424 N$22848 N$22847 "Straight Waveguide" sch_x=-207 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11425 N$22850 N$22849 "Straight Waveguide" sch_x=-207 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11426 N$22852 N$22851 "Straight Waveguide" sch_x=-207 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11427 N$22854 N$22853 "Straight Waveguide" sch_x=-207 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11428 N$22856 N$22855 "Straight Waveguide" sch_x=-207 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11429 N$22858 N$22857 "Straight Waveguide" sch_x=-207 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11430 N$22860 N$22859 "Straight Waveguide" sch_x=-207 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11431 N$22862 N$22861 "Straight Waveguide" sch_x=-207 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11432 N$22864 N$22863 "Straight Waveguide" sch_x=-207 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11433 N$22866 N$22865 "Straight Waveguide" sch_x=-205 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11434 N$22868 N$22867 "Straight Waveguide" sch_x=-205 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11435 N$22870 N$22869 "Straight Waveguide" sch_x=-205 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11436 N$22872 N$22871 "Straight Waveguide" sch_x=-205 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11437 N$22874 N$22873 "Straight Waveguide" sch_x=-205 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11438 N$22876 N$22875 "Straight Waveguide" sch_x=-205 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11439 N$22878 N$22877 "Straight Waveguide" sch_x=-205 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11440 N$22880 N$22879 "Straight Waveguide" sch_x=-205 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11441 N$22882 N$22881 "Straight Waveguide" sch_x=-205 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11442 N$22884 N$22883 "Straight Waveguide" sch_x=-205 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11443 N$22886 N$22885 "Straight Waveguide" sch_x=-205 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11444 N$22888 N$22887 "Straight Waveguide" sch_x=-205 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11445 N$22890 N$22889 "Straight Waveguide" sch_x=-205 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11446 N$22892 N$22891 "Straight Waveguide" sch_x=-205 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11447 N$22894 N$22893 "Straight Waveguide" sch_x=-205 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11448 N$22896 N$22895 "Straight Waveguide" sch_x=-205 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11449 N$22898 N$22897 "Straight Waveguide" sch_x=-205 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11450 N$22900 N$22899 "Straight Waveguide" sch_x=-205 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11451 N$22902 N$22901 "Straight Waveguide" sch_x=-205 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11452 N$22904 N$22903 "Straight Waveguide" sch_x=-205 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11453 N$22906 N$22905 "Straight Waveguide" sch_x=-205 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11454 N$22908 N$22907 "Straight Waveguide" sch_x=-205 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11455 N$22910 N$22909 "Straight Waveguide" sch_x=-205 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11456 N$22912 N$22911 "Straight Waveguide" sch_x=-205 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11457 N$22914 N$22913 "Straight Waveguide" sch_x=-205 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11458 N$22916 N$22915 "Straight Waveguide" sch_x=-205 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11459 N$22918 N$22917 "Straight Waveguide" sch_x=-205 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11460 N$22920 N$22919 "Straight Waveguide" sch_x=-205 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11461 N$22922 N$22921 "Straight Waveguide" sch_x=-205 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11462 N$22924 N$22923 "Straight Waveguide" sch_x=-205 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11463 N$22926 N$22925 "Straight Waveguide" sch_x=-205 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11464 N$22928 N$22927 "Straight Waveguide" sch_x=-205 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11465 N$22930 N$22929 "Straight Waveguide" sch_x=-205 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11466 N$22932 N$22931 "Straight Waveguide" sch_x=-205 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11467 N$22934 N$22933 "Straight Waveguide" sch_x=-205 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11468 N$22936 N$22935 "Straight Waveguide" sch_x=-205 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11469 N$22938 N$22937 "Straight Waveguide" sch_x=-205 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11470 N$22940 N$22939 "Straight Waveguide" sch_x=-205 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11471 N$22942 N$22941 "Straight Waveguide" sch_x=-205 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11472 N$22944 N$22943 "Straight Waveguide" sch_x=-205 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11473 N$22946 N$22945 "Straight Waveguide" sch_x=-205 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11474 N$22948 N$22947 "Straight Waveguide" sch_x=-205 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11475 N$22950 N$22949 "Straight Waveguide" sch_x=-205 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11476 N$22952 N$22951 "Straight Waveguide" sch_x=-205 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11477 N$22954 N$22953 "Straight Waveguide" sch_x=-205 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11478 N$22956 N$22955 "Straight Waveguide" sch_x=-205 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11479 N$22958 N$22957 "Straight Waveguide" sch_x=-205 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11480 N$22960 N$22959 "Straight Waveguide" sch_x=-205 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11481 N$22962 N$22961 "Straight Waveguide" sch_x=-205 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11482 N$22964 N$22963 "Straight Waveguide" sch_x=-205 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11483 N$22966 N$22965 "Straight Waveguide" sch_x=-205 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11484 N$22968 N$22967 "Straight Waveguide" sch_x=-205 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11485 N$22970 N$22969 "Straight Waveguide" sch_x=-205 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11486 N$22972 N$22971 "Straight Waveguide" sch_x=-205 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11487 N$22974 N$22973 "Straight Waveguide" sch_x=-205 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11488 N$22976 N$22975 "Straight Waveguide" sch_x=-205 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11489 N$22978 N$22977 "Straight Waveguide" sch_x=-205 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11490 N$22980 N$22979 "Straight Waveguide" sch_x=-205 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11491 N$22982 N$22981 "Straight Waveguide" sch_x=-205 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11492 N$22984 N$22983 "Straight Waveguide" sch_x=-205 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11493 N$22986 N$22985 "Straight Waveguide" sch_x=-205 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11494 N$22988 N$22987 "Straight Waveguide" sch_x=-205 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11495 N$22990 N$22989 "Straight Waveguide" sch_x=-205 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11496 N$22992 N$22991 "Straight Waveguide" sch_x=-205 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11497 N$22994 N$22993 "Straight Waveguide" sch_x=-205 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11498 N$22996 N$22995 "Straight Waveguide" sch_x=-205 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11499 N$22998 N$22997 "Straight Waveguide" sch_x=-205 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11500 N$23000 N$22999 "Straight Waveguide" sch_x=-205 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11501 N$23002 N$23001 "Straight Waveguide" sch_x=-205 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11502 N$23004 N$23003 "Straight Waveguide" sch_x=-205 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11503 N$23006 N$23005 "Straight Waveguide" sch_x=-205 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11504 N$23008 N$23007 "Straight Waveguide" sch_x=-205 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11505 N$23010 N$23009 "Straight Waveguide" sch_x=-205 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11506 N$23012 N$23011 "Straight Waveguide" sch_x=-205 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11507 N$23014 N$23013 "Straight Waveguide" sch_x=-205 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11508 N$23016 N$23015 "Straight Waveguide" sch_x=-205 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11509 N$23018 N$23017 "Straight Waveguide" sch_x=-205 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11510 N$23020 N$23019 "Straight Waveguide" sch_x=-205 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11511 N$23022 N$23021 "Straight Waveguide" sch_x=-203 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11512 N$23024 N$23023 "Straight Waveguide" sch_x=-203 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11513 N$23026 N$23025 "Straight Waveguide" sch_x=-203 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11514 N$23028 N$23027 "Straight Waveguide" sch_x=-203 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11515 N$23030 N$23029 "Straight Waveguide" sch_x=-203 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11516 N$23032 N$23031 "Straight Waveguide" sch_x=-203 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11517 N$23034 N$23033 "Straight Waveguide" sch_x=-203 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11518 N$23036 N$23035 "Straight Waveguide" sch_x=-203 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11519 N$23038 N$23037 "Straight Waveguide" sch_x=-203 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11520 N$23040 N$23039 "Straight Waveguide" sch_x=-203 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11521 N$23042 N$23041 "Straight Waveguide" sch_x=-203 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11522 N$23044 N$23043 "Straight Waveguide" sch_x=-203 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11523 N$23046 N$23045 "Straight Waveguide" sch_x=-203 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11524 N$23048 N$23047 "Straight Waveguide" sch_x=-203 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11525 N$23050 N$23049 "Straight Waveguide" sch_x=-203 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11526 N$23052 N$23051 "Straight Waveguide" sch_x=-203 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11527 N$23054 N$23053 "Straight Waveguide" sch_x=-203 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11528 N$23056 N$23055 "Straight Waveguide" sch_x=-203 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11529 N$23058 N$23057 "Straight Waveguide" sch_x=-203 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11530 N$23060 N$23059 "Straight Waveguide" sch_x=-203 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11531 N$23062 N$23061 "Straight Waveguide" sch_x=-203 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11532 N$23064 N$23063 "Straight Waveguide" sch_x=-203 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11533 N$23066 N$23065 "Straight Waveguide" sch_x=-203 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11534 N$23068 N$23067 "Straight Waveguide" sch_x=-203 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11535 N$23070 N$23069 "Straight Waveguide" sch_x=-203 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11536 N$23072 N$23071 "Straight Waveguide" sch_x=-203 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11537 N$23074 N$23073 "Straight Waveguide" sch_x=-203 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11538 N$23076 N$23075 "Straight Waveguide" sch_x=-203 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11539 N$23078 N$23077 "Straight Waveguide" sch_x=-203 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11540 N$23080 N$23079 "Straight Waveguide" sch_x=-203 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11541 N$23082 N$23081 "Straight Waveguide" sch_x=-203 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11542 N$23084 N$23083 "Straight Waveguide" sch_x=-203 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11543 N$23086 N$23085 "Straight Waveguide" sch_x=-203 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11544 N$23088 N$23087 "Straight Waveguide" sch_x=-203 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11545 N$23090 N$23089 "Straight Waveguide" sch_x=-203 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11546 N$23092 N$23091 "Straight Waveguide" sch_x=-203 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11547 N$23094 N$23093 "Straight Waveguide" sch_x=-203 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11548 N$23096 N$23095 "Straight Waveguide" sch_x=-203 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11549 N$23098 N$23097 "Straight Waveguide" sch_x=-203 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11550 N$23100 N$23099 "Straight Waveguide" sch_x=-203 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11551 N$23102 N$23101 "Straight Waveguide" sch_x=-203 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11552 N$23104 N$23103 "Straight Waveguide" sch_x=-203 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11553 N$23106 N$23105 "Straight Waveguide" sch_x=-203 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11554 N$23108 N$23107 "Straight Waveguide" sch_x=-203 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11555 N$23110 N$23109 "Straight Waveguide" sch_x=-203 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11556 N$23112 N$23111 "Straight Waveguide" sch_x=-203 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11557 N$23114 N$23113 "Straight Waveguide" sch_x=-203 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11558 N$23116 N$23115 "Straight Waveguide" sch_x=-203 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11559 N$23118 N$23117 "Straight Waveguide" sch_x=-203 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11560 N$23120 N$23119 "Straight Waveguide" sch_x=-203 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11561 N$23122 N$23121 "Straight Waveguide" sch_x=-203 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11562 N$23124 N$23123 "Straight Waveguide" sch_x=-203 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11563 N$23126 N$23125 "Straight Waveguide" sch_x=-203 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11564 N$23128 N$23127 "Straight Waveguide" sch_x=-203 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11565 N$23130 N$23129 "Straight Waveguide" sch_x=-203 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11566 N$23132 N$23131 "Straight Waveguide" sch_x=-203 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11567 N$23134 N$23133 "Straight Waveguide" sch_x=-203 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11568 N$23136 N$23135 "Straight Waveguide" sch_x=-203 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11569 N$23138 N$23137 "Straight Waveguide" sch_x=-203 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11570 N$23140 N$23139 "Straight Waveguide" sch_x=-203 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11571 N$23142 N$23141 "Straight Waveguide" sch_x=-203 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11572 N$23144 N$23143 "Straight Waveguide" sch_x=-203 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11573 N$23146 N$23145 "Straight Waveguide" sch_x=-203 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11574 N$23148 N$23147 "Straight Waveguide" sch_x=-203 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11575 N$23150 N$23149 "Straight Waveguide" sch_x=-203 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11576 N$23152 N$23151 "Straight Waveguide" sch_x=-203 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11577 N$23154 N$23153 "Straight Waveguide" sch_x=-203 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11578 N$23156 N$23155 "Straight Waveguide" sch_x=-203 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11579 N$23158 N$23157 "Straight Waveguide" sch_x=-203 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11580 N$23160 N$23159 "Straight Waveguide" sch_x=-203 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11581 N$23162 N$23161 "Straight Waveguide" sch_x=-203 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11582 N$23164 N$23163 "Straight Waveguide" sch_x=-203 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11583 N$23166 N$23165 "Straight Waveguide" sch_x=-203 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11584 N$23168 N$23167 "Straight Waveguide" sch_x=-203 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11585 N$23170 N$23169 "Straight Waveguide" sch_x=-203 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11586 N$23172 N$23171 "Straight Waveguide" sch_x=-203 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11587 N$23174 N$23173 "Straight Waveguide" sch_x=-201 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11588 N$23176 N$23175 "Straight Waveguide" sch_x=-201 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11589 N$23178 N$23177 "Straight Waveguide" sch_x=-201 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11590 N$23180 N$23179 "Straight Waveguide" sch_x=-201 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11591 N$23182 N$23181 "Straight Waveguide" sch_x=-201 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11592 N$23184 N$23183 "Straight Waveguide" sch_x=-201 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11593 N$23186 N$23185 "Straight Waveguide" sch_x=-201 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11594 N$23188 N$23187 "Straight Waveguide" sch_x=-201 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11595 N$23190 N$23189 "Straight Waveguide" sch_x=-201 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11596 N$23192 N$23191 "Straight Waveguide" sch_x=-201 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11597 N$23194 N$23193 "Straight Waveguide" sch_x=-201 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11598 N$23196 N$23195 "Straight Waveguide" sch_x=-201 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11599 N$23198 N$23197 "Straight Waveguide" sch_x=-201 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11600 N$23200 N$23199 "Straight Waveguide" sch_x=-201 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11601 N$23202 N$23201 "Straight Waveguide" sch_x=-201 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11602 N$23204 N$23203 "Straight Waveguide" sch_x=-201 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11603 N$23206 N$23205 "Straight Waveguide" sch_x=-201 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11604 N$23208 N$23207 "Straight Waveguide" sch_x=-201 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11605 N$23210 N$23209 "Straight Waveguide" sch_x=-201 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11606 N$23212 N$23211 "Straight Waveguide" sch_x=-201 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11607 N$23214 N$23213 "Straight Waveguide" sch_x=-201 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11608 N$23216 N$23215 "Straight Waveguide" sch_x=-201 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11609 N$23218 N$23217 "Straight Waveguide" sch_x=-201 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11610 N$23220 N$23219 "Straight Waveguide" sch_x=-201 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11611 N$23222 N$23221 "Straight Waveguide" sch_x=-201 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11612 N$23224 N$23223 "Straight Waveguide" sch_x=-201 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11613 N$23226 N$23225 "Straight Waveguide" sch_x=-201 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11614 N$23228 N$23227 "Straight Waveguide" sch_x=-201 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11615 N$23230 N$23229 "Straight Waveguide" sch_x=-201 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11616 N$23232 N$23231 "Straight Waveguide" sch_x=-201 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11617 N$23234 N$23233 "Straight Waveguide" sch_x=-201 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11618 N$23236 N$23235 "Straight Waveguide" sch_x=-201 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11619 N$23238 N$23237 "Straight Waveguide" sch_x=-201 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11620 N$23240 N$23239 "Straight Waveguide" sch_x=-201 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11621 N$23242 N$23241 "Straight Waveguide" sch_x=-201 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11622 N$23244 N$23243 "Straight Waveguide" sch_x=-201 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11623 N$23246 N$23245 "Straight Waveguide" sch_x=-201 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11624 N$23248 N$23247 "Straight Waveguide" sch_x=-201 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11625 N$23250 N$23249 "Straight Waveguide" sch_x=-201 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11626 N$23252 N$23251 "Straight Waveguide" sch_x=-201 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11627 N$23254 N$23253 "Straight Waveguide" sch_x=-201 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11628 N$23256 N$23255 "Straight Waveguide" sch_x=-201 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11629 N$23258 N$23257 "Straight Waveguide" sch_x=-201 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11630 N$23260 N$23259 "Straight Waveguide" sch_x=-201 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11631 N$23262 N$23261 "Straight Waveguide" sch_x=-201 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11632 N$23264 N$23263 "Straight Waveguide" sch_x=-201 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11633 N$23266 N$23265 "Straight Waveguide" sch_x=-201 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11634 N$23268 N$23267 "Straight Waveguide" sch_x=-201 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11635 N$23270 N$23269 "Straight Waveguide" sch_x=-201 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11636 N$23272 N$23271 "Straight Waveguide" sch_x=-201 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11637 N$23274 N$23273 "Straight Waveguide" sch_x=-201 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11638 N$23276 N$23275 "Straight Waveguide" sch_x=-201 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11639 N$23278 N$23277 "Straight Waveguide" sch_x=-201 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11640 N$23280 N$23279 "Straight Waveguide" sch_x=-201 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11641 N$23282 N$23281 "Straight Waveguide" sch_x=-201 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11642 N$23284 N$23283 "Straight Waveguide" sch_x=-201 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11643 N$23286 N$23285 "Straight Waveguide" sch_x=-201 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11644 N$23288 N$23287 "Straight Waveguide" sch_x=-201 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11645 N$23290 N$23289 "Straight Waveguide" sch_x=-201 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11646 N$23292 N$23291 "Straight Waveguide" sch_x=-201 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11647 N$23294 N$23293 "Straight Waveguide" sch_x=-201 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11648 N$23296 N$23295 "Straight Waveguide" sch_x=-201 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11649 N$23298 N$23297 "Straight Waveguide" sch_x=-201 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11650 N$23300 N$23299 "Straight Waveguide" sch_x=-201 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11651 N$23302 N$23301 "Straight Waveguide" sch_x=-201 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11652 N$23304 N$23303 "Straight Waveguide" sch_x=-201 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11653 N$23306 N$23305 "Straight Waveguide" sch_x=-201 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11654 N$23308 N$23307 "Straight Waveguide" sch_x=-201 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11655 N$23310 N$23309 "Straight Waveguide" sch_x=-201 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11656 N$23312 N$23311 "Straight Waveguide" sch_x=-201 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11657 N$23314 N$23313 "Straight Waveguide" sch_x=-201 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11658 N$23316 N$23315 "Straight Waveguide" sch_x=-201 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11659 N$23318 N$23317 "Straight Waveguide" sch_x=-201 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11660 N$23320 N$23319 "Straight Waveguide" sch_x=-201 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11661 N$23322 N$23321 "Straight Waveguide" sch_x=-199 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11662 N$23324 N$23323 "Straight Waveguide" sch_x=-199 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11663 N$23326 N$23325 "Straight Waveguide" sch_x=-199 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11664 N$23328 N$23327 "Straight Waveguide" sch_x=-199 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11665 N$23330 N$23329 "Straight Waveguide" sch_x=-199 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11666 N$23332 N$23331 "Straight Waveguide" sch_x=-199 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11667 N$23334 N$23333 "Straight Waveguide" sch_x=-199 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11668 N$23336 N$23335 "Straight Waveguide" sch_x=-199 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11669 N$23338 N$23337 "Straight Waveguide" sch_x=-199 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11670 N$23340 N$23339 "Straight Waveguide" sch_x=-199 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11671 N$23342 N$23341 "Straight Waveguide" sch_x=-199 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11672 N$23344 N$23343 "Straight Waveguide" sch_x=-199 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11673 N$23346 N$23345 "Straight Waveguide" sch_x=-199 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11674 N$23348 N$23347 "Straight Waveguide" sch_x=-199 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11675 N$23350 N$23349 "Straight Waveguide" sch_x=-199 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11676 N$23352 N$23351 "Straight Waveguide" sch_x=-199 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11677 N$23354 N$23353 "Straight Waveguide" sch_x=-199 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11678 N$23356 N$23355 "Straight Waveguide" sch_x=-199 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11679 N$23358 N$23357 "Straight Waveguide" sch_x=-199 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11680 N$23360 N$23359 "Straight Waveguide" sch_x=-199 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11681 N$23362 N$23361 "Straight Waveguide" sch_x=-199 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11682 N$23364 N$23363 "Straight Waveguide" sch_x=-199 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11683 N$23366 N$23365 "Straight Waveguide" sch_x=-199 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11684 N$23368 N$23367 "Straight Waveguide" sch_x=-199 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11685 N$23370 N$23369 "Straight Waveguide" sch_x=-199 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11686 N$23372 N$23371 "Straight Waveguide" sch_x=-199 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11687 N$23374 N$23373 "Straight Waveguide" sch_x=-199 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11688 N$23376 N$23375 "Straight Waveguide" sch_x=-199 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11689 N$23378 N$23377 "Straight Waveguide" sch_x=-199 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11690 N$23380 N$23379 "Straight Waveguide" sch_x=-199 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11691 N$23382 N$23381 "Straight Waveguide" sch_x=-199 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11692 N$23384 N$23383 "Straight Waveguide" sch_x=-199 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11693 N$23386 N$23385 "Straight Waveguide" sch_x=-199 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11694 N$23388 N$23387 "Straight Waveguide" sch_x=-199 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11695 N$23390 N$23389 "Straight Waveguide" sch_x=-199 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11696 N$23392 N$23391 "Straight Waveguide" sch_x=-199 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11697 N$23394 N$23393 "Straight Waveguide" sch_x=-199 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11698 N$23396 N$23395 "Straight Waveguide" sch_x=-199 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11699 N$23398 N$23397 "Straight Waveguide" sch_x=-199 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11700 N$23400 N$23399 "Straight Waveguide" sch_x=-199 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11701 N$23402 N$23401 "Straight Waveguide" sch_x=-199 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11702 N$23404 N$23403 "Straight Waveguide" sch_x=-199 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11703 N$23406 N$23405 "Straight Waveguide" sch_x=-199 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11704 N$23408 N$23407 "Straight Waveguide" sch_x=-199 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11705 N$23410 N$23409 "Straight Waveguide" sch_x=-199 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11706 N$23412 N$23411 "Straight Waveguide" sch_x=-199 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11707 N$23414 N$23413 "Straight Waveguide" sch_x=-199 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11708 N$23416 N$23415 "Straight Waveguide" sch_x=-199 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11709 N$23418 N$23417 "Straight Waveguide" sch_x=-199 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11710 N$23420 N$23419 "Straight Waveguide" sch_x=-199 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11711 N$23422 N$23421 "Straight Waveguide" sch_x=-199 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11712 N$23424 N$23423 "Straight Waveguide" sch_x=-199 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11713 N$23426 N$23425 "Straight Waveguide" sch_x=-199 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11714 N$23428 N$23427 "Straight Waveguide" sch_x=-199 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11715 N$23430 N$23429 "Straight Waveguide" sch_x=-199 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11716 N$23432 N$23431 "Straight Waveguide" sch_x=-199 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11717 N$23434 N$23433 "Straight Waveguide" sch_x=-199 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11718 N$23436 N$23435 "Straight Waveguide" sch_x=-199 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11719 N$23438 N$23437 "Straight Waveguide" sch_x=-199 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11720 N$23440 N$23439 "Straight Waveguide" sch_x=-199 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11721 N$23442 N$23441 "Straight Waveguide" sch_x=-199 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11722 N$23444 N$23443 "Straight Waveguide" sch_x=-199 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11723 N$23446 N$23445 "Straight Waveguide" sch_x=-199 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11724 N$23448 N$23447 "Straight Waveguide" sch_x=-199 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11725 N$23450 N$23449 "Straight Waveguide" sch_x=-199 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11726 N$23452 N$23451 "Straight Waveguide" sch_x=-199 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11727 N$23454 N$23453 "Straight Waveguide" sch_x=-199 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11728 N$23456 N$23455 "Straight Waveguide" sch_x=-199 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11729 N$23458 N$23457 "Straight Waveguide" sch_x=-199 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11730 N$23460 N$23459 "Straight Waveguide" sch_x=-199 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11731 N$23462 N$23461 "Straight Waveguide" sch_x=-199 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11732 N$23464 N$23463 "Straight Waveguide" sch_x=-199 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11733 N$23466 N$23465 "Straight Waveguide" sch_x=-197 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11734 N$23468 N$23467 "Straight Waveguide" sch_x=-197 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11735 N$23470 N$23469 "Straight Waveguide" sch_x=-197 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11736 N$23472 N$23471 "Straight Waveguide" sch_x=-197 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11737 N$23474 N$23473 "Straight Waveguide" sch_x=-197 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11738 N$23476 N$23475 "Straight Waveguide" sch_x=-197 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11739 N$23478 N$23477 "Straight Waveguide" sch_x=-197 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11740 N$23480 N$23479 "Straight Waveguide" sch_x=-197 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11741 N$23482 N$23481 "Straight Waveguide" sch_x=-197 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11742 N$23484 N$23483 "Straight Waveguide" sch_x=-197 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11743 N$23486 N$23485 "Straight Waveguide" sch_x=-197 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11744 N$23488 N$23487 "Straight Waveguide" sch_x=-197 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11745 N$23490 N$23489 "Straight Waveguide" sch_x=-197 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11746 N$23492 N$23491 "Straight Waveguide" sch_x=-197 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11747 N$23494 N$23493 "Straight Waveguide" sch_x=-197 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11748 N$23496 N$23495 "Straight Waveguide" sch_x=-197 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11749 N$23498 N$23497 "Straight Waveguide" sch_x=-197 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11750 N$23500 N$23499 "Straight Waveguide" sch_x=-197 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11751 N$23502 N$23501 "Straight Waveguide" sch_x=-197 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11752 N$23504 N$23503 "Straight Waveguide" sch_x=-197 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11753 N$23506 N$23505 "Straight Waveguide" sch_x=-197 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11754 N$23508 N$23507 "Straight Waveguide" sch_x=-197 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11755 N$23510 N$23509 "Straight Waveguide" sch_x=-197 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11756 N$23512 N$23511 "Straight Waveguide" sch_x=-197 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11757 N$23514 N$23513 "Straight Waveguide" sch_x=-197 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11758 N$23516 N$23515 "Straight Waveguide" sch_x=-197 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11759 N$23518 N$23517 "Straight Waveguide" sch_x=-197 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11760 N$23520 N$23519 "Straight Waveguide" sch_x=-197 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11761 N$23522 N$23521 "Straight Waveguide" sch_x=-197 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11762 N$23524 N$23523 "Straight Waveguide" sch_x=-197 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11763 N$23526 N$23525 "Straight Waveguide" sch_x=-197 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11764 N$23528 N$23527 "Straight Waveguide" sch_x=-197 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11765 N$23530 N$23529 "Straight Waveguide" sch_x=-197 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11766 N$23532 N$23531 "Straight Waveguide" sch_x=-197 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11767 N$23534 N$23533 "Straight Waveguide" sch_x=-197 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11768 N$23536 N$23535 "Straight Waveguide" sch_x=-197 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11769 N$23538 N$23537 "Straight Waveguide" sch_x=-197 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11770 N$23540 N$23539 "Straight Waveguide" sch_x=-197 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11771 N$23542 N$23541 "Straight Waveguide" sch_x=-197 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11772 N$23544 N$23543 "Straight Waveguide" sch_x=-197 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11773 N$23546 N$23545 "Straight Waveguide" sch_x=-197 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11774 N$23548 N$23547 "Straight Waveguide" sch_x=-197 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11775 N$23550 N$23549 "Straight Waveguide" sch_x=-197 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11776 N$23552 N$23551 "Straight Waveguide" sch_x=-197 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11777 N$23554 N$23553 "Straight Waveguide" sch_x=-197 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11778 N$23556 N$23555 "Straight Waveguide" sch_x=-197 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11779 N$23558 N$23557 "Straight Waveguide" sch_x=-197 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11780 N$23560 N$23559 "Straight Waveguide" sch_x=-197 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11781 N$23562 N$23561 "Straight Waveguide" sch_x=-197 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11782 N$23564 N$23563 "Straight Waveguide" sch_x=-197 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11783 N$23566 N$23565 "Straight Waveguide" sch_x=-197 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11784 N$23568 N$23567 "Straight Waveguide" sch_x=-197 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11785 N$23570 N$23569 "Straight Waveguide" sch_x=-197 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11786 N$23572 N$23571 "Straight Waveguide" sch_x=-197 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11787 N$23574 N$23573 "Straight Waveguide" sch_x=-197 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11788 N$23576 N$23575 "Straight Waveguide" sch_x=-197 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11789 N$23578 N$23577 "Straight Waveguide" sch_x=-197 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11790 N$23580 N$23579 "Straight Waveguide" sch_x=-197 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11791 N$23582 N$23581 "Straight Waveguide" sch_x=-197 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11792 N$23584 N$23583 "Straight Waveguide" sch_x=-197 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11793 N$23586 N$23585 "Straight Waveguide" sch_x=-197 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11794 N$23588 N$23587 "Straight Waveguide" sch_x=-197 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11795 N$23590 N$23589 "Straight Waveguide" sch_x=-197 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11796 N$23592 N$23591 "Straight Waveguide" sch_x=-197 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11797 N$23594 N$23593 "Straight Waveguide" sch_x=-197 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11798 N$23596 N$23595 "Straight Waveguide" sch_x=-197 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11799 N$23598 N$23597 "Straight Waveguide" sch_x=-197 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11800 N$23600 N$23599 "Straight Waveguide" sch_x=-197 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11801 N$23602 N$23601 "Straight Waveguide" sch_x=-197 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11802 N$23604 N$23603 "Straight Waveguide" sch_x=-197 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11803 N$23606 N$23605 "Straight Waveguide" sch_x=-195 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11804 N$23608 N$23607 "Straight Waveguide" sch_x=-195 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11805 N$23610 N$23609 "Straight Waveguide" sch_x=-195 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11806 N$23612 N$23611 "Straight Waveguide" sch_x=-195 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11807 N$23614 N$23613 "Straight Waveguide" sch_x=-195 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11808 N$23616 N$23615 "Straight Waveguide" sch_x=-195 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11809 N$23618 N$23617 "Straight Waveguide" sch_x=-195 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11810 N$23620 N$23619 "Straight Waveguide" sch_x=-195 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11811 N$23622 N$23621 "Straight Waveguide" sch_x=-195 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11812 N$23624 N$23623 "Straight Waveguide" sch_x=-195 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11813 N$23626 N$23625 "Straight Waveguide" sch_x=-195 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11814 N$23628 N$23627 "Straight Waveguide" sch_x=-195 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11815 N$23630 N$23629 "Straight Waveguide" sch_x=-195 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11816 N$23632 N$23631 "Straight Waveguide" sch_x=-195 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11817 N$23634 N$23633 "Straight Waveguide" sch_x=-195 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11818 N$23636 N$23635 "Straight Waveguide" sch_x=-195 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11819 N$23638 N$23637 "Straight Waveguide" sch_x=-195 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11820 N$23640 N$23639 "Straight Waveguide" sch_x=-195 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11821 N$23642 N$23641 "Straight Waveguide" sch_x=-195 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11822 N$23644 N$23643 "Straight Waveguide" sch_x=-195 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11823 N$23646 N$23645 "Straight Waveguide" sch_x=-195 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11824 N$23648 N$23647 "Straight Waveguide" sch_x=-195 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11825 N$23650 N$23649 "Straight Waveguide" sch_x=-195 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11826 N$23652 N$23651 "Straight Waveguide" sch_x=-195 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11827 N$23654 N$23653 "Straight Waveguide" sch_x=-195 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11828 N$23656 N$23655 "Straight Waveguide" sch_x=-195 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11829 N$23658 N$23657 "Straight Waveguide" sch_x=-195 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11830 N$23660 N$23659 "Straight Waveguide" sch_x=-195 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11831 N$23662 N$23661 "Straight Waveguide" sch_x=-195 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11832 N$23664 N$23663 "Straight Waveguide" sch_x=-195 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11833 N$23666 N$23665 "Straight Waveguide" sch_x=-195 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11834 N$23668 N$23667 "Straight Waveguide" sch_x=-195 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11835 N$23670 N$23669 "Straight Waveguide" sch_x=-195 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11836 N$23672 N$23671 "Straight Waveguide" sch_x=-195 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11837 N$23674 N$23673 "Straight Waveguide" sch_x=-195 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11838 N$23676 N$23675 "Straight Waveguide" sch_x=-195 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11839 N$23678 N$23677 "Straight Waveguide" sch_x=-195 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11840 N$23680 N$23679 "Straight Waveguide" sch_x=-195 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11841 N$23682 N$23681 "Straight Waveguide" sch_x=-195 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11842 N$23684 N$23683 "Straight Waveguide" sch_x=-195 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11843 N$23686 N$23685 "Straight Waveguide" sch_x=-195 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11844 N$23688 N$23687 "Straight Waveguide" sch_x=-195 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11845 N$23690 N$23689 "Straight Waveguide" sch_x=-195 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11846 N$23692 N$23691 "Straight Waveguide" sch_x=-195 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11847 N$23694 N$23693 "Straight Waveguide" sch_x=-195 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11848 N$23696 N$23695 "Straight Waveguide" sch_x=-195 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11849 N$23698 N$23697 "Straight Waveguide" sch_x=-195 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11850 N$23700 N$23699 "Straight Waveguide" sch_x=-195 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11851 N$23702 N$23701 "Straight Waveguide" sch_x=-195 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11852 N$23704 N$23703 "Straight Waveguide" sch_x=-195 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11853 N$23706 N$23705 "Straight Waveguide" sch_x=-195 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11854 N$23708 N$23707 "Straight Waveguide" sch_x=-195 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11855 N$23710 N$23709 "Straight Waveguide" sch_x=-195 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11856 N$23712 N$23711 "Straight Waveguide" sch_x=-195 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11857 N$23714 N$23713 "Straight Waveguide" sch_x=-195 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11858 N$23716 N$23715 "Straight Waveguide" sch_x=-195 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11859 N$23718 N$23717 "Straight Waveguide" sch_x=-195 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11860 N$23720 N$23719 "Straight Waveguide" sch_x=-195 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11861 N$23722 N$23721 "Straight Waveguide" sch_x=-195 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11862 N$23724 N$23723 "Straight Waveguide" sch_x=-195 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11863 N$23726 N$23725 "Straight Waveguide" sch_x=-195 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11864 N$23728 N$23727 "Straight Waveguide" sch_x=-195 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11865 N$23730 N$23729 "Straight Waveguide" sch_x=-195 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11866 N$23732 N$23731 "Straight Waveguide" sch_x=-195 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11867 N$23734 N$23733 "Straight Waveguide" sch_x=-195 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11868 N$23736 N$23735 "Straight Waveguide" sch_x=-195 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11869 N$23738 N$23737 "Straight Waveguide" sch_x=-195 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11870 N$23740 N$23739 "Straight Waveguide" sch_x=-195 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11871 N$23742 N$23741 "Straight Waveguide" sch_x=-193 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11872 N$23744 N$23743 "Straight Waveguide" sch_x=-193 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11873 N$23746 N$23745 "Straight Waveguide" sch_x=-193 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11874 N$23748 N$23747 "Straight Waveguide" sch_x=-193 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11875 N$23750 N$23749 "Straight Waveguide" sch_x=-193 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11876 N$23752 N$23751 "Straight Waveguide" sch_x=-193 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11877 N$23754 N$23753 "Straight Waveguide" sch_x=-193 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11878 N$23756 N$23755 "Straight Waveguide" sch_x=-193 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11879 N$23758 N$23757 "Straight Waveguide" sch_x=-193 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11880 N$23760 N$23759 "Straight Waveguide" sch_x=-193 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11881 N$23762 N$23761 "Straight Waveguide" sch_x=-193 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11882 N$23764 N$23763 "Straight Waveguide" sch_x=-193 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11883 N$23766 N$23765 "Straight Waveguide" sch_x=-193 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11884 N$23768 N$23767 "Straight Waveguide" sch_x=-193 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11885 N$23770 N$23769 "Straight Waveguide" sch_x=-193 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11886 N$23772 N$23771 "Straight Waveguide" sch_x=-193 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11887 N$23774 N$23773 "Straight Waveguide" sch_x=-193 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11888 N$23776 N$23775 "Straight Waveguide" sch_x=-193 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11889 N$23778 N$23777 "Straight Waveguide" sch_x=-193 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11890 N$23780 N$23779 "Straight Waveguide" sch_x=-193 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11891 N$23782 N$23781 "Straight Waveguide" sch_x=-193 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11892 N$23784 N$23783 "Straight Waveguide" sch_x=-193 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11893 N$23786 N$23785 "Straight Waveguide" sch_x=-193 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11894 N$23788 N$23787 "Straight Waveguide" sch_x=-193 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11895 N$23790 N$23789 "Straight Waveguide" sch_x=-193 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11896 N$23792 N$23791 "Straight Waveguide" sch_x=-193 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11897 N$23794 N$23793 "Straight Waveguide" sch_x=-193 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11898 N$23796 N$23795 "Straight Waveguide" sch_x=-193 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11899 N$23798 N$23797 "Straight Waveguide" sch_x=-193 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11900 N$23800 N$23799 "Straight Waveguide" sch_x=-193 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11901 N$23802 N$23801 "Straight Waveguide" sch_x=-193 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11902 N$23804 N$23803 "Straight Waveguide" sch_x=-193 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11903 N$23806 N$23805 "Straight Waveguide" sch_x=-193 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11904 N$23808 N$23807 "Straight Waveguide" sch_x=-193 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11905 N$23810 N$23809 "Straight Waveguide" sch_x=-193 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11906 N$23812 N$23811 "Straight Waveguide" sch_x=-193 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11907 N$23814 N$23813 "Straight Waveguide" sch_x=-193 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11908 N$23816 N$23815 "Straight Waveguide" sch_x=-193 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11909 N$23818 N$23817 "Straight Waveguide" sch_x=-193 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11910 N$23820 N$23819 "Straight Waveguide" sch_x=-193 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11911 N$23822 N$23821 "Straight Waveguide" sch_x=-193 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11912 N$23824 N$23823 "Straight Waveguide" sch_x=-193 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11913 N$23826 N$23825 "Straight Waveguide" sch_x=-193 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11914 N$23828 N$23827 "Straight Waveguide" sch_x=-193 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11915 N$23830 N$23829 "Straight Waveguide" sch_x=-193 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11916 N$23832 N$23831 "Straight Waveguide" sch_x=-193 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11917 N$23834 N$23833 "Straight Waveguide" sch_x=-193 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11918 N$23836 N$23835 "Straight Waveguide" sch_x=-193 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11919 N$23838 N$23837 "Straight Waveguide" sch_x=-193 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11920 N$23840 N$23839 "Straight Waveguide" sch_x=-193 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11921 N$23842 N$23841 "Straight Waveguide" sch_x=-193 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11922 N$23844 N$23843 "Straight Waveguide" sch_x=-193 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11923 N$23846 N$23845 "Straight Waveguide" sch_x=-193 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11924 N$23848 N$23847 "Straight Waveguide" sch_x=-193 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11925 N$23850 N$23849 "Straight Waveguide" sch_x=-193 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11926 N$23852 N$23851 "Straight Waveguide" sch_x=-193 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11927 N$23854 N$23853 "Straight Waveguide" sch_x=-193 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11928 N$23856 N$23855 "Straight Waveguide" sch_x=-193 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11929 N$23858 N$23857 "Straight Waveguide" sch_x=-193 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11930 N$23860 N$23859 "Straight Waveguide" sch_x=-193 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11931 N$23862 N$23861 "Straight Waveguide" sch_x=-193 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11932 N$23864 N$23863 "Straight Waveguide" sch_x=-193 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11933 N$23866 N$23865 "Straight Waveguide" sch_x=-193 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11934 N$23868 N$23867 "Straight Waveguide" sch_x=-193 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11935 N$23870 N$23869 "Straight Waveguide" sch_x=-193 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11936 N$23872 N$23871 "Straight Waveguide" sch_x=-193 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11937 N$23874 N$23873 "Straight Waveguide" sch_x=-191 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11938 N$23876 N$23875 "Straight Waveguide" sch_x=-191 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11939 N$23878 N$23877 "Straight Waveguide" sch_x=-191 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11940 N$23880 N$23879 "Straight Waveguide" sch_x=-191 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11941 N$23882 N$23881 "Straight Waveguide" sch_x=-191 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11942 N$23884 N$23883 "Straight Waveguide" sch_x=-191 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11943 N$23886 N$23885 "Straight Waveguide" sch_x=-191 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11944 N$23888 N$23887 "Straight Waveguide" sch_x=-191 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11945 N$23890 N$23889 "Straight Waveguide" sch_x=-191 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11946 N$23892 N$23891 "Straight Waveguide" sch_x=-191 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11947 N$23894 N$23893 "Straight Waveguide" sch_x=-191 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11948 N$23896 N$23895 "Straight Waveguide" sch_x=-191 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11949 N$23898 N$23897 "Straight Waveguide" sch_x=-191 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11950 N$23900 N$23899 "Straight Waveguide" sch_x=-191 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11951 N$23902 N$23901 "Straight Waveguide" sch_x=-191 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11952 N$23904 N$23903 "Straight Waveguide" sch_x=-191 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11953 N$23906 N$23905 "Straight Waveguide" sch_x=-191 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11954 N$23908 N$23907 "Straight Waveguide" sch_x=-191 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11955 N$23910 N$23909 "Straight Waveguide" sch_x=-191 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11956 N$23912 N$23911 "Straight Waveguide" sch_x=-191 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11957 N$23914 N$23913 "Straight Waveguide" sch_x=-191 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11958 N$23916 N$23915 "Straight Waveguide" sch_x=-191 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11959 N$23918 N$23917 "Straight Waveguide" sch_x=-191 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11960 N$23920 N$23919 "Straight Waveguide" sch_x=-191 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11961 N$23922 N$23921 "Straight Waveguide" sch_x=-191 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11962 N$23924 N$23923 "Straight Waveguide" sch_x=-191 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11963 N$23926 N$23925 "Straight Waveguide" sch_x=-191 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11964 N$23928 N$23927 "Straight Waveguide" sch_x=-191 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11965 N$23930 N$23929 "Straight Waveguide" sch_x=-191 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11966 N$23932 N$23931 "Straight Waveguide" sch_x=-191 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11967 N$23934 N$23933 "Straight Waveguide" sch_x=-191 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11968 N$23936 N$23935 "Straight Waveguide" sch_x=-191 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11969 N$23938 N$23937 "Straight Waveguide" sch_x=-191 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11970 N$23940 N$23939 "Straight Waveguide" sch_x=-191 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11971 N$23942 N$23941 "Straight Waveguide" sch_x=-191 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11972 N$23944 N$23943 "Straight Waveguide" sch_x=-191 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11973 N$23946 N$23945 "Straight Waveguide" sch_x=-191 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11974 N$23948 N$23947 "Straight Waveguide" sch_x=-191 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11975 N$23950 N$23949 "Straight Waveguide" sch_x=-191 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11976 N$23952 N$23951 "Straight Waveguide" sch_x=-191 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11977 N$23954 N$23953 "Straight Waveguide" sch_x=-191 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11978 N$23956 N$23955 "Straight Waveguide" sch_x=-191 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11979 N$23958 N$23957 "Straight Waveguide" sch_x=-191 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11980 N$23960 N$23959 "Straight Waveguide" sch_x=-191 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11981 N$23962 N$23961 "Straight Waveguide" sch_x=-191 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11982 N$23964 N$23963 "Straight Waveguide" sch_x=-191 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11983 N$23966 N$23965 "Straight Waveguide" sch_x=-191 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11984 N$23968 N$23967 "Straight Waveguide" sch_x=-191 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11985 N$23970 N$23969 "Straight Waveguide" sch_x=-191 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11986 N$23972 N$23971 "Straight Waveguide" sch_x=-191 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11987 N$23974 N$23973 "Straight Waveguide" sch_x=-191 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11988 N$23976 N$23975 "Straight Waveguide" sch_x=-191 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11989 N$23978 N$23977 "Straight Waveguide" sch_x=-191 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11990 N$23980 N$23979 "Straight Waveguide" sch_x=-191 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11991 N$23982 N$23981 "Straight Waveguide" sch_x=-191 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11992 N$23984 N$23983 "Straight Waveguide" sch_x=-191 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11993 N$23986 N$23985 "Straight Waveguide" sch_x=-191 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11994 N$23988 N$23987 "Straight Waveguide" sch_x=-191 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11995 N$23990 N$23989 "Straight Waveguide" sch_x=-191 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11996 N$23992 N$23991 "Straight Waveguide" sch_x=-191 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11997 N$23994 N$23993 "Straight Waveguide" sch_x=-191 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11998 N$23996 N$23995 "Straight Waveguide" sch_x=-191 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11999 N$23998 N$23997 "Straight Waveguide" sch_x=-191 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12000 N$24000 N$23999 "Straight Waveguide" sch_x=-191 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12001 N$24002 N$24001 "Straight Waveguide" sch_x=-189 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12002 N$24004 N$24003 "Straight Waveguide" sch_x=-189 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12003 N$24006 N$24005 "Straight Waveguide" sch_x=-189 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12004 N$24008 N$24007 "Straight Waveguide" sch_x=-189 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12005 N$24010 N$24009 "Straight Waveguide" sch_x=-189 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12006 N$24012 N$24011 "Straight Waveguide" sch_x=-189 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12007 N$24014 N$24013 "Straight Waveguide" sch_x=-189 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12008 N$24016 N$24015 "Straight Waveguide" sch_x=-189 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12009 N$24018 N$24017 "Straight Waveguide" sch_x=-189 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12010 N$24020 N$24019 "Straight Waveguide" sch_x=-189 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12011 N$24022 N$24021 "Straight Waveguide" sch_x=-189 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12012 N$24024 N$24023 "Straight Waveguide" sch_x=-189 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12013 N$24026 N$24025 "Straight Waveguide" sch_x=-189 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12014 N$24028 N$24027 "Straight Waveguide" sch_x=-189 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12015 N$24030 N$24029 "Straight Waveguide" sch_x=-189 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12016 N$24032 N$24031 "Straight Waveguide" sch_x=-189 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12017 N$24034 N$24033 "Straight Waveguide" sch_x=-189 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12018 N$24036 N$24035 "Straight Waveguide" sch_x=-189 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12019 N$24038 N$24037 "Straight Waveguide" sch_x=-189 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12020 N$24040 N$24039 "Straight Waveguide" sch_x=-189 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12021 N$24042 N$24041 "Straight Waveguide" sch_x=-189 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12022 N$24044 N$24043 "Straight Waveguide" sch_x=-189 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12023 N$24046 N$24045 "Straight Waveguide" sch_x=-189 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12024 N$24048 N$24047 "Straight Waveguide" sch_x=-189 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12025 N$24050 N$24049 "Straight Waveguide" sch_x=-189 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12026 N$24052 N$24051 "Straight Waveguide" sch_x=-189 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12027 N$24054 N$24053 "Straight Waveguide" sch_x=-189 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12028 N$24056 N$24055 "Straight Waveguide" sch_x=-189 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12029 N$24058 N$24057 "Straight Waveguide" sch_x=-189 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12030 N$24060 N$24059 "Straight Waveguide" sch_x=-189 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12031 N$24062 N$24061 "Straight Waveguide" sch_x=-189 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12032 N$24064 N$24063 "Straight Waveguide" sch_x=-189 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12033 N$24066 N$24065 "Straight Waveguide" sch_x=-189 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12034 N$24068 N$24067 "Straight Waveguide" sch_x=-189 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12035 N$24070 N$24069 "Straight Waveguide" sch_x=-189 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12036 N$24072 N$24071 "Straight Waveguide" sch_x=-189 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12037 N$24074 N$24073 "Straight Waveguide" sch_x=-189 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12038 N$24076 N$24075 "Straight Waveguide" sch_x=-189 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12039 N$24078 N$24077 "Straight Waveguide" sch_x=-189 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12040 N$24080 N$24079 "Straight Waveguide" sch_x=-189 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12041 N$24082 N$24081 "Straight Waveguide" sch_x=-189 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12042 N$24084 N$24083 "Straight Waveguide" sch_x=-189 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12043 N$24086 N$24085 "Straight Waveguide" sch_x=-189 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12044 N$24088 N$24087 "Straight Waveguide" sch_x=-189 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12045 N$24090 N$24089 "Straight Waveguide" sch_x=-189 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12046 N$24092 N$24091 "Straight Waveguide" sch_x=-189 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12047 N$24094 N$24093 "Straight Waveguide" sch_x=-189 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12048 N$24096 N$24095 "Straight Waveguide" sch_x=-189 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12049 N$24098 N$24097 "Straight Waveguide" sch_x=-189 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12050 N$24100 N$24099 "Straight Waveguide" sch_x=-189 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12051 N$24102 N$24101 "Straight Waveguide" sch_x=-189 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12052 N$24104 N$24103 "Straight Waveguide" sch_x=-189 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12053 N$24106 N$24105 "Straight Waveguide" sch_x=-189 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12054 N$24108 N$24107 "Straight Waveguide" sch_x=-189 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12055 N$24110 N$24109 "Straight Waveguide" sch_x=-189 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12056 N$24112 N$24111 "Straight Waveguide" sch_x=-189 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12057 N$24114 N$24113 "Straight Waveguide" sch_x=-189 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12058 N$24116 N$24115 "Straight Waveguide" sch_x=-189 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12059 N$24118 N$24117 "Straight Waveguide" sch_x=-189 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12060 N$24120 N$24119 "Straight Waveguide" sch_x=-189 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12061 N$24122 N$24121 "Straight Waveguide" sch_x=-189 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12062 N$24124 N$24123 "Straight Waveguide" sch_x=-189 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12063 N$24126 N$24125 "Straight Waveguide" sch_x=-187 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12064 N$24128 N$24127 "Straight Waveguide" sch_x=-187 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12065 N$24130 N$24129 "Straight Waveguide" sch_x=-187 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12066 N$24132 N$24131 "Straight Waveguide" sch_x=-187 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12067 N$24134 N$24133 "Straight Waveguide" sch_x=-187 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12068 N$24136 N$24135 "Straight Waveguide" sch_x=-187 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12069 N$24138 N$24137 "Straight Waveguide" sch_x=-187 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12070 N$24140 N$24139 "Straight Waveguide" sch_x=-187 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12071 N$24142 N$24141 "Straight Waveguide" sch_x=-187 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12072 N$24144 N$24143 "Straight Waveguide" sch_x=-187 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12073 N$24146 N$24145 "Straight Waveguide" sch_x=-187 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12074 N$24148 N$24147 "Straight Waveguide" sch_x=-187 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12075 N$24150 N$24149 "Straight Waveguide" sch_x=-187 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12076 N$24152 N$24151 "Straight Waveguide" sch_x=-187 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12077 N$24154 N$24153 "Straight Waveguide" sch_x=-187 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12078 N$24156 N$24155 "Straight Waveguide" sch_x=-187 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12079 N$24158 N$24157 "Straight Waveguide" sch_x=-187 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12080 N$24160 N$24159 "Straight Waveguide" sch_x=-187 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12081 N$24162 N$24161 "Straight Waveguide" sch_x=-187 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12082 N$24164 N$24163 "Straight Waveguide" sch_x=-187 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12083 N$24166 N$24165 "Straight Waveguide" sch_x=-187 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12084 N$24168 N$24167 "Straight Waveguide" sch_x=-187 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12085 N$24170 N$24169 "Straight Waveguide" sch_x=-187 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12086 N$24172 N$24171 "Straight Waveguide" sch_x=-187 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12087 N$24174 N$24173 "Straight Waveguide" sch_x=-187 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12088 N$24176 N$24175 "Straight Waveguide" sch_x=-187 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12089 N$24178 N$24177 "Straight Waveguide" sch_x=-187 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12090 N$24180 N$24179 "Straight Waveguide" sch_x=-187 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12091 N$24182 N$24181 "Straight Waveguide" sch_x=-187 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12092 N$24184 N$24183 "Straight Waveguide" sch_x=-187 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12093 N$24186 N$24185 "Straight Waveguide" sch_x=-187 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12094 N$24188 N$24187 "Straight Waveguide" sch_x=-187 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12095 N$24190 N$24189 "Straight Waveguide" sch_x=-187 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12096 N$24192 N$24191 "Straight Waveguide" sch_x=-187 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12097 N$24194 N$24193 "Straight Waveguide" sch_x=-187 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12098 N$24196 N$24195 "Straight Waveguide" sch_x=-187 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12099 N$24198 N$24197 "Straight Waveguide" sch_x=-187 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12100 N$24200 N$24199 "Straight Waveguide" sch_x=-187 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12101 N$24202 N$24201 "Straight Waveguide" sch_x=-187 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12102 N$24204 N$24203 "Straight Waveguide" sch_x=-187 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12103 N$24206 N$24205 "Straight Waveguide" sch_x=-187 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12104 N$24208 N$24207 "Straight Waveguide" sch_x=-187 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12105 N$24210 N$24209 "Straight Waveguide" sch_x=-187 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12106 N$24212 N$24211 "Straight Waveguide" sch_x=-187 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12107 N$24214 N$24213 "Straight Waveguide" sch_x=-187 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12108 N$24216 N$24215 "Straight Waveguide" sch_x=-187 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12109 N$24218 N$24217 "Straight Waveguide" sch_x=-187 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12110 N$24220 N$24219 "Straight Waveguide" sch_x=-187 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12111 N$24222 N$24221 "Straight Waveguide" sch_x=-187 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12112 N$24224 N$24223 "Straight Waveguide" sch_x=-187 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12113 N$24226 N$24225 "Straight Waveguide" sch_x=-187 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12114 N$24228 N$24227 "Straight Waveguide" sch_x=-187 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12115 N$24230 N$24229 "Straight Waveguide" sch_x=-187 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12116 N$24232 N$24231 "Straight Waveguide" sch_x=-187 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12117 N$24234 N$24233 "Straight Waveguide" sch_x=-187 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12118 N$24236 N$24235 "Straight Waveguide" sch_x=-187 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12119 N$24238 N$24237 "Straight Waveguide" sch_x=-187 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12120 N$24240 N$24239 "Straight Waveguide" sch_x=-187 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12121 N$24242 N$24241 "Straight Waveguide" sch_x=-187 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12122 N$24244 N$24243 "Straight Waveguide" sch_x=-187 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12123 N$24246 N$24245 "Straight Waveguide" sch_x=-185 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12124 N$24248 N$24247 "Straight Waveguide" sch_x=-185 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12125 N$24250 N$24249 "Straight Waveguide" sch_x=-185 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12126 N$24252 N$24251 "Straight Waveguide" sch_x=-185 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12127 N$24254 N$24253 "Straight Waveguide" sch_x=-185 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12128 N$24256 N$24255 "Straight Waveguide" sch_x=-185 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12129 N$24258 N$24257 "Straight Waveguide" sch_x=-185 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12130 N$24260 N$24259 "Straight Waveguide" sch_x=-185 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12131 N$24262 N$24261 "Straight Waveguide" sch_x=-185 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12132 N$24264 N$24263 "Straight Waveguide" sch_x=-185 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12133 N$24266 N$24265 "Straight Waveguide" sch_x=-185 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12134 N$24268 N$24267 "Straight Waveguide" sch_x=-185 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12135 N$24270 N$24269 "Straight Waveguide" sch_x=-185 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12136 N$24272 N$24271 "Straight Waveguide" sch_x=-185 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12137 N$24274 N$24273 "Straight Waveguide" sch_x=-185 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12138 N$24276 N$24275 "Straight Waveguide" sch_x=-185 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12139 N$24278 N$24277 "Straight Waveguide" sch_x=-185 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12140 N$24280 N$24279 "Straight Waveguide" sch_x=-185 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12141 N$24282 N$24281 "Straight Waveguide" sch_x=-185 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12142 N$24284 N$24283 "Straight Waveguide" sch_x=-185 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12143 N$24286 N$24285 "Straight Waveguide" sch_x=-185 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12144 N$24288 N$24287 "Straight Waveguide" sch_x=-185 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12145 N$24290 N$24289 "Straight Waveguide" sch_x=-185 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12146 N$24292 N$24291 "Straight Waveguide" sch_x=-185 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12147 N$24294 N$24293 "Straight Waveguide" sch_x=-185 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12148 N$24296 N$24295 "Straight Waveguide" sch_x=-185 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12149 N$24298 N$24297 "Straight Waveguide" sch_x=-185 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12150 N$24300 N$24299 "Straight Waveguide" sch_x=-185 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12151 N$24302 N$24301 "Straight Waveguide" sch_x=-185 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12152 N$24304 N$24303 "Straight Waveguide" sch_x=-185 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12153 N$24306 N$24305 "Straight Waveguide" sch_x=-185 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12154 N$24308 N$24307 "Straight Waveguide" sch_x=-185 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12155 N$24310 N$24309 "Straight Waveguide" sch_x=-185 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12156 N$24312 N$24311 "Straight Waveguide" sch_x=-185 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12157 N$24314 N$24313 "Straight Waveguide" sch_x=-185 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12158 N$24316 N$24315 "Straight Waveguide" sch_x=-185 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12159 N$24318 N$24317 "Straight Waveguide" sch_x=-185 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12160 N$24320 N$24319 "Straight Waveguide" sch_x=-185 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12161 N$24322 N$24321 "Straight Waveguide" sch_x=-185 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12162 N$24324 N$24323 "Straight Waveguide" sch_x=-185 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12163 N$24326 N$24325 "Straight Waveguide" sch_x=-185 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12164 N$24328 N$24327 "Straight Waveguide" sch_x=-185 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12165 N$24330 N$24329 "Straight Waveguide" sch_x=-185 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12166 N$24332 N$24331 "Straight Waveguide" sch_x=-185 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12167 N$24334 N$24333 "Straight Waveguide" sch_x=-185 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12168 N$24336 N$24335 "Straight Waveguide" sch_x=-185 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12169 N$24338 N$24337 "Straight Waveguide" sch_x=-185 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12170 N$24340 N$24339 "Straight Waveguide" sch_x=-185 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12171 N$24342 N$24341 "Straight Waveguide" sch_x=-185 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12172 N$24344 N$24343 "Straight Waveguide" sch_x=-185 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12173 N$24346 N$24345 "Straight Waveguide" sch_x=-185 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12174 N$24348 N$24347 "Straight Waveguide" sch_x=-185 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12175 N$24350 N$24349 "Straight Waveguide" sch_x=-185 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12176 N$24352 N$24351 "Straight Waveguide" sch_x=-185 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12177 N$24354 N$24353 "Straight Waveguide" sch_x=-185 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12178 N$24356 N$24355 "Straight Waveguide" sch_x=-185 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12179 N$24358 N$24357 "Straight Waveguide" sch_x=-185 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12180 N$24360 N$24359 "Straight Waveguide" sch_x=-185 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12181 N$24362 N$24361 "Straight Waveguide" sch_x=-183 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12182 N$24364 N$24363 "Straight Waveguide" sch_x=-183 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12183 N$24366 N$24365 "Straight Waveguide" sch_x=-183 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12184 N$24368 N$24367 "Straight Waveguide" sch_x=-183 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12185 N$24370 N$24369 "Straight Waveguide" sch_x=-183 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12186 N$24372 N$24371 "Straight Waveguide" sch_x=-183 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12187 N$24374 N$24373 "Straight Waveguide" sch_x=-183 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12188 N$24376 N$24375 "Straight Waveguide" sch_x=-183 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12189 N$24378 N$24377 "Straight Waveguide" sch_x=-183 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12190 N$24380 N$24379 "Straight Waveguide" sch_x=-183 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12191 N$24382 N$24381 "Straight Waveguide" sch_x=-183 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12192 N$24384 N$24383 "Straight Waveguide" sch_x=-183 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12193 N$24386 N$24385 "Straight Waveguide" sch_x=-183 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12194 N$24388 N$24387 "Straight Waveguide" sch_x=-183 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12195 N$24390 N$24389 "Straight Waveguide" sch_x=-183 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12196 N$24392 N$24391 "Straight Waveguide" sch_x=-183 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12197 N$24394 N$24393 "Straight Waveguide" sch_x=-183 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12198 N$24396 N$24395 "Straight Waveguide" sch_x=-183 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12199 N$24398 N$24397 "Straight Waveguide" sch_x=-183 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12200 N$24400 N$24399 "Straight Waveguide" sch_x=-183 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12201 N$24402 N$24401 "Straight Waveguide" sch_x=-183 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12202 N$24404 N$24403 "Straight Waveguide" sch_x=-183 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12203 N$24406 N$24405 "Straight Waveguide" sch_x=-183 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12204 N$24408 N$24407 "Straight Waveguide" sch_x=-183 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12205 N$24410 N$24409 "Straight Waveguide" sch_x=-183 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12206 N$24412 N$24411 "Straight Waveguide" sch_x=-183 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12207 N$24414 N$24413 "Straight Waveguide" sch_x=-183 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12208 N$24416 N$24415 "Straight Waveguide" sch_x=-183 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12209 N$24418 N$24417 "Straight Waveguide" sch_x=-183 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12210 N$24420 N$24419 "Straight Waveguide" sch_x=-183 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12211 N$24422 N$24421 "Straight Waveguide" sch_x=-183 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12212 N$24424 N$24423 "Straight Waveguide" sch_x=-183 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12213 N$24426 N$24425 "Straight Waveguide" sch_x=-183 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12214 N$24428 N$24427 "Straight Waveguide" sch_x=-183 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12215 N$24430 N$24429 "Straight Waveguide" sch_x=-183 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12216 N$24432 N$24431 "Straight Waveguide" sch_x=-183 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12217 N$24434 N$24433 "Straight Waveguide" sch_x=-183 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12218 N$24436 N$24435 "Straight Waveguide" sch_x=-183 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12219 N$24438 N$24437 "Straight Waveguide" sch_x=-183 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12220 N$24440 N$24439 "Straight Waveguide" sch_x=-183 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12221 N$24442 N$24441 "Straight Waveguide" sch_x=-183 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12222 N$24444 N$24443 "Straight Waveguide" sch_x=-183 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12223 N$24446 N$24445 "Straight Waveguide" sch_x=-183 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12224 N$24448 N$24447 "Straight Waveguide" sch_x=-183 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12225 N$24450 N$24449 "Straight Waveguide" sch_x=-183 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12226 N$24452 N$24451 "Straight Waveguide" sch_x=-183 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12227 N$24454 N$24453 "Straight Waveguide" sch_x=-183 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12228 N$24456 N$24455 "Straight Waveguide" sch_x=-183 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12229 N$24458 N$24457 "Straight Waveguide" sch_x=-183 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12230 N$24460 N$24459 "Straight Waveguide" sch_x=-183 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12231 N$24462 N$24461 "Straight Waveguide" sch_x=-183 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12232 N$24464 N$24463 "Straight Waveguide" sch_x=-183 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12233 N$24466 N$24465 "Straight Waveguide" sch_x=-183 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12234 N$24468 N$24467 "Straight Waveguide" sch_x=-183 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12235 N$24470 N$24469 "Straight Waveguide" sch_x=-183 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12236 N$24472 N$24471 "Straight Waveguide" sch_x=-183 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12237 N$24474 N$24473 "Straight Waveguide" sch_x=-181 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12238 N$24476 N$24475 "Straight Waveguide" sch_x=-181 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12239 N$24478 N$24477 "Straight Waveguide" sch_x=-181 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12240 N$24480 N$24479 "Straight Waveguide" sch_x=-181 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12241 N$24482 N$24481 "Straight Waveguide" sch_x=-181 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12242 N$24484 N$24483 "Straight Waveguide" sch_x=-181 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12243 N$24486 N$24485 "Straight Waveguide" sch_x=-181 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12244 N$24488 N$24487 "Straight Waveguide" sch_x=-181 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12245 N$24490 N$24489 "Straight Waveguide" sch_x=-181 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12246 N$24492 N$24491 "Straight Waveguide" sch_x=-181 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12247 N$24494 N$24493 "Straight Waveguide" sch_x=-181 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12248 N$24496 N$24495 "Straight Waveguide" sch_x=-181 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12249 N$24498 N$24497 "Straight Waveguide" sch_x=-181 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12250 N$24500 N$24499 "Straight Waveguide" sch_x=-181 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12251 N$24502 N$24501 "Straight Waveguide" sch_x=-181 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12252 N$24504 N$24503 "Straight Waveguide" sch_x=-181 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12253 N$24506 N$24505 "Straight Waveguide" sch_x=-181 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12254 N$24508 N$24507 "Straight Waveguide" sch_x=-181 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12255 N$24510 N$24509 "Straight Waveguide" sch_x=-181 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12256 N$24512 N$24511 "Straight Waveguide" sch_x=-181 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12257 N$24514 N$24513 "Straight Waveguide" sch_x=-181 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12258 N$24516 N$24515 "Straight Waveguide" sch_x=-181 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12259 N$24518 N$24517 "Straight Waveguide" sch_x=-181 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12260 N$24520 N$24519 "Straight Waveguide" sch_x=-181 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12261 N$24522 N$24521 "Straight Waveguide" sch_x=-181 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12262 N$24524 N$24523 "Straight Waveguide" sch_x=-181 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12263 N$24526 N$24525 "Straight Waveguide" sch_x=-181 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12264 N$24528 N$24527 "Straight Waveguide" sch_x=-181 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12265 N$24530 N$24529 "Straight Waveguide" sch_x=-181 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12266 N$24532 N$24531 "Straight Waveguide" sch_x=-181 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12267 N$24534 N$24533 "Straight Waveguide" sch_x=-181 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12268 N$24536 N$24535 "Straight Waveguide" sch_x=-181 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12269 N$24538 N$24537 "Straight Waveguide" sch_x=-181 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12270 N$24540 N$24539 "Straight Waveguide" sch_x=-181 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12271 N$24542 N$24541 "Straight Waveguide" sch_x=-181 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12272 N$24544 N$24543 "Straight Waveguide" sch_x=-181 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12273 N$24546 N$24545 "Straight Waveguide" sch_x=-181 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12274 N$24548 N$24547 "Straight Waveguide" sch_x=-181 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12275 N$24550 N$24549 "Straight Waveguide" sch_x=-181 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12276 N$24552 N$24551 "Straight Waveguide" sch_x=-181 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12277 N$24554 N$24553 "Straight Waveguide" sch_x=-181 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12278 N$24556 N$24555 "Straight Waveguide" sch_x=-181 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12279 N$24558 N$24557 "Straight Waveguide" sch_x=-181 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12280 N$24560 N$24559 "Straight Waveguide" sch_x=-181 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12281 N$24562 N$24561 "Straight Waveguide" sch_x=-181 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12282 N$24564 N$24563 "Straight Waveguide" sch_x=-181 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12283 N$24566 N$24565 "Straight Waveguide" sch_x=-181 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12284 N$24568 N$24567 "Straight Waveguide" sch_x=-181 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12285 N$24570 N$24569 "Straight Waveguide" sch_x=-181 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12286 N$24572 N$24571 "Straight Waveguide" sch_x=-181 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12287 N$24574 N$24573 "Straight Waveguide" sch_x=-181 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12288 N$24576 N$24575 "Straight Waveguide" sch_x=-181 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12289 N$24578 N$24577 "Straight Waveguide" sch_x=-181 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12290 N$24580 N$24579 "Straight Waveguide" sch_x=-181 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12291 N$24582 N$24581 "Straight Waveguide" sch_x=-179 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12292 N$24584 N$24583 "Straight Waveguide" sch_x=-179 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12293 N$24586 N$24585 "Straight Waveguide" sch_x=-179 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12294 N$24588 N$24587 "Straight Waveguide" sch_x=-179 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12295 N$24590 N$24589 "Straight Waveguide" sch_x=-179 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12296 N$24592 N$24591 "Straight Waveguide" sch_x=-179 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12297 N$24594 N$24593 "Straight Waveguide" sch_x=-179 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12298 N$24596 N$24595 "Straight Waveguide" sch_x=-179 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12299 N$24598 N$24597 "Straight Waveguide" sch_x=-179 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12300 N$24600 N$24599 "Straight Waveguide" sch_x=-179 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12301 N$24602 N$24601 "Straight Waveguide" sch_x=-179 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12302 N$24604 N$24603 "Straight Waveguide" sch_x=-179 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12303 N$24606 N$24605 "Straight Waveguide" sch_x=-179 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12304 N$24608 N$24607 "Straight Waveguide" sch_x=-179 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12305 N$24610 N$24609 "Straight Waveguide" sch_x=-179 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12306 N$24612 N$24611 "Straight Waveguide" sch_x=-179 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12307 N$24614 N$24613 "Straight Waveguide" sch_x=-179 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12308 N$24616 N$24615 "Straight Waveguide" sch_x=-179 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12309 N$24618 N$24617 "Straight Waveguide" sch_x=-179 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12310 N$24620 N$24619 "Straight Waveguide" sch_x=-179 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12311 N$24622 N$24621 "Straight Waveguide" sch_x=-179 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12312 N$24624 N$24623 "Straight Waveguide" sch_x=-179 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12313 N$24626 N$24625 "Straight Waveguide" sch_x=-179 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12314 N$24628 N$24627 "Straight Waveguide" sch_x=-179 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12315 N$24630 N$24629 "Straight Waveguide" sch_x=-179 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12316 N$24632 N$24631 "Straight Waveguide" sch_x=-179 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12317 N$24634 N$24633 "Straight Waveguide" sch_x=-179 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12318 N$24636 N$24635 "Straight Waveguide" sch_x=-179 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12319 N$24638 N$24637 "Straight Waveguide" sch_x=-179 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12320 N$24640 N$24639 "Straight Waveguide" sch_x=-179 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12321 N$24642 N$24641 "Straight Waveguide" sch_x=-179 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12322 N$24644 N$24643 "Straight Waveguide" sch_x=-179 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12323 N$24646 N$24645 "Straight Waveguide" sch_x=-179 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12324 N$24648 N$24647 "Straight Waveguide" sch_x=-179 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12325 N$24650 N$24649 "Straight Waveguide" sch_x=-179 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12326 N$24652 N$24651 "Straight Waveguide" sch_x=-179 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12327 N$24654 N$24653 "Straight Waveguide" sch_x=-179 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12328 N$24656 N$24655 "Straight Waveguide" sch_x=-179 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12329 N$24658 N$24657 "Straight Waveguide" sch_x=-179 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12330 N$24660 N$24659 "Straight Waveguide" sch_x=-179 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12331 N$24662 N$24661 "Straight Waveguide" sch_x=-179 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12332 N$24664 N$24663 "Straight Waveguide" sch_x=-179 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12333 N$24666 N$24665 "Straight Waveguide" sch_x=-179 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12334 N$24668 N$24667 "Straight Waveguide" sch_x=-179 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12335 N$24670 N$24669 "Straight Waveguide" sch_x=-179 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12336 N$24672 N$24671 "Straight Waveguide" sch_x=-179 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12337 N$24674 N$24673 "Straight Waveguide" sch_x=-179 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12338 N$24676 N$24675 "Straight Waveguide" sch_x=-179 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12339 N$24678 N$24677 "Straight Waveguide" sch_x=-179 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12340 N$24680 N$24679 "Straight Waveguide" sch_x=-179 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12341 N$24682 N$24681 "Straight Waveguide" sch_x=-179 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12342 N$24684 N$24683 "Straight Waveguide" sch_x=-179 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12343 N$24686 N$24685 "Straight Waveguide" sch_x=-177 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12344 N$24688 N$24687 "Straight Waveguide" sch_x=-177 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12345 N$24690 N$24689 "Straight Waveguide" sch_x=-177 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12346 N$24692 N$24691 "Straight Waveguide" sch_x=-177 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12347 N$24694 N$24693 "Straight Waveguide" sch_x=-177 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12348 N$24696 N$24695 "Straight Waveguide" sch_x=-177 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12349 N$24698 N$24697 "Straight Waveguide" sch_x=-177 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12350 N$24700 N$24699 "Straight Waveguide" sch_x=-177 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12351 N$24702 N$24701 "Straight Waveguide" sch_x=-177 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12352 N$24704 N$24703 "Straight Waveguide" sch_x=-177 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12353 N$24706 N$24705 "Straight Waveguide" sch_x=-177 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12354 N$24708 N$24707 "Straight Waveguide" sch_x=-177 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12355 N$24710 N$24709 "Straight Waveguide" sch_x=-177 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12356 N$24712 N$24711 "Straight Waveguide" sch_x=-177 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12357 N$24714 N$24713 "Straight Waveguide" sch_x=-177 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12358 N$24716 N$24715 "Straight Waveguide" sch_x=-177 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12359 N$24718 N$24717 "Straight Waveguide" sch_x=-177 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12360 N$24720 N$24719 "Straight Waveguide" sch_x=-177 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12361 N$24722 N$24721 "Straight Waveguide" sch_x=-177 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12362 N$24724 N$24723 "Straight Waveguide" sch_x=-177 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12363 N$24726 N$24725 "Straight Waveguide" sch_x=-177 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12364 N$24728 N$24727 "Straight Waveguide" sch_x=-177 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12365 N$24730 N$24729 "Straight Waveguide" sch_x=-177 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12366 N$24732 N$24731 "Straight Waveguide" sch_x=-177 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12367 N$24734 N$24733 "Straight Waveguide" sch_x=-177 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12368 N$24736 N$24735 "Straight Waveguide" sch_x=-177 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12369 N$24738 N$24737 "Straight Waveguide" sch_x=-177 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12370 N$24740 N$24739 "Straight Waveguide" sch_x=-177 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12371 N$24742 N$24741 "Straight Waveguide" sch_x=-177 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12372 N$24744 N$24743 "Straight Waveguide" sch_x=-177 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12373 N$24746 N$24745 "Straight Waveguide" sch_x=-177 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12374 N$24748 N$24747 "Straight Waveguide" sch_x=-177 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12375 N$24750 N$24749 "Straight Waveguide" sch_x=-177 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12376 N$24752 N$24751 "Straight Waveguide" sch_x=-177 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12377 N$24754 N$24753 "Straight Waveguide" sch_x=-177 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12378 N$24756 N$24755 "Straight Waveguide" sch_x=-177 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12379 N$24758 N$24757 "Straight Waveguide" sch_x=-177 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12380 N$24760 N$24759 "Straight Waveguide" sch_x=-177 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12381 N$24762 N$24761 "Straight Waveguide" sch_x=-177 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12382 N$24764 N$24763 "Straight Waveguide" sch_x=-177 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12383 N$24766 N$24765 "Straight Waveguide" sch_x=-177 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12384 N$24768 N$24767 "Straight Waveguide" sch_x=-177 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12385 N$24770 N$24769 "Straight Waveguide" sch_x=-177 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12386 N$24772 N$24771 "Straight Waveguide" sch_x=-177 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12387 N$24774 N$24773 "Straight Waveguide" sch_x=-177 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12388 N$24776 N$24775 "Straight Waveguide" sch_x=-177 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12389 N$24778 N$24777 "Straight Waveguide" sch_x=-177 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12390 N$24780 N$24779 "Straight Waveguide" sch_x=-177 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12391 N$24782 N$24781 "Straight Waveguide" sch_x=-177 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12392 N$24784 N$24783 "Straight Waveguide" sch_x=-177 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12393 N$24786 N$24785 "Straight Waveguide" sch_x=-175 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12394 N$24788 N$24787 "Straight Waveguide" sch_x=-175 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12395 N$24790 N$24789 "Straight Waveguide" sch_x=-175 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12396 N$24792 N$24791 "Straight Waveguide" sch_x=-175 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12397 N$24794 N$24793 "Straight Waveguide" sch_x=-175 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12398 N$24796 N$24795 "Straight Waveguide" sch_x=-175 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12399 N$24798 N$24797 "Straight Waveguide" sch_x=-175 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12400 N$24800 N$24799 "Straight Waveguide" sch_x=-175 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12401 N$24802 N$24801 "Straight Waveguide" sch_x=-175 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12402 N$24804 N$24803 "Straight Waveguide" sch_x=-175 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12403 N$24806 N$24805 "Straight Waveguide" sch_x=-175 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12404 N$24808 N$24807 "Straight Waveguide" sch_x=-175 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12405 N$24810 N$24809 "Straight Waveguide" sch_x=-175 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12406 N$24812 N$24811 "Straight Waveguide" sch_x=-175 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12407 N$24814 N$24813 "Straight Waveguide" sch_x=-175 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12408 N$24816 N$24815 "Straight Waveguide" sch_x=-175 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12409 N$24818 N$24817 "Straight Waveguide" sch_x=-175 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12410 N$24820 N$24819 "Straight Waveguide" sch_x=-175 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12411 N$24822 N$24821 "Straight Waveguide" sch_x=-175 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12412 N$24824 N$24823 "Straight Waveguide" sch_x=-175 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12413 N$24826 N$24825 "Straight Waveguide" sch_x=-175 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12414 N$24828 N$24827 "Straight Waveguide" sch_x=-175 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12415 N$24830 N$24829 "Straight Waveguide" sch_x=-175 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12416 N$24832 N$24831 "Straight Waveguide" sch_x=-175 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12417 N$24834 N$24833 "Straight Waveguide" sch_x=-175 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12418 N$24836 N$24835 "Straight Waveguide" sch_x=-175 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12419 N$24838 N$24837 "Straight Waveguide" sch_x=-175 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12420 N$24840 N$24839 "Straight Waveguide" sch_x=-175 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12421 N$24842 N$24841 "Straight Waveguide" sch_x=-175 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12422 N$24844 N$24843 "Straight Waveguide" sch_x=-175 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12423 N$24846 N$24845 "Straight Waveguide" sch_x=-175 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12424 N$24848 N$24847 "Straight Waveguide" sch_x=-175 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12425 N$24850 N$24849 "Straight Waveguide" sch_x=-175 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12426 N$24852 N$24851 "Straight Waveguide" sch_x=-175 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12427 N$24854 N$24853 "Straight Waveguide" sch_x=-175 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12428 N$24856 N$24855 "Straight Waveguide" sch_x=-175 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12429 N$24858 N$24857 "Straight Waveguide" sch_x=-175 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12430 N$24860 N$24859 "Straight Waveguide" sch_x=-175 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12431 N$24862 N$24861 "Straight Waveguide" sch_x=-175 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12432 N$24864 N$24863 "Straight Waveguide" sch_x=-175 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12433 N$24866 N$24865 "Straight Waveguide" sch_x=-175 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12434 N$24868 N$24867 "Straight Waveguide" sch_x=-175 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12435 N$24870 N$24869 "Straight Waveguide" sch_x=-175 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12436 N$24872 N$24871 "Straight Waveguide" sch_x=-175 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12437 N$24874 N$24873 "Straight Waveguide" sch_x=-175 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12438 N$24876 N$24875 "Straight Waveguide" sch_x=-175 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12439 N$24878 N$24877 "Straight Waveguide" sch_x=-175 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12440 N$24880 N$24879 "Straight Waveguide" sch_x=-175 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12441 N$24882 N$24881 "Straight Waveguide" sch_x=-173 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12442 N$24884 N$24883 "Straight Waveguide" sch_x=-173 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12443 N$24886 N$24885 "Straight Waveguide" sch_x=-173 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12444 N$24888 N$24887 "Straight Waveguide" sch_x=-173 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12445 N$24890 N$24889 "Straight Waveguide" sch_x=-173 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12446 N$24892 N$24891 "Straight Waveguide" sch_x=-173 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12447 N$24894 N$24893 "Straight Waveguide" sch_x=-173 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12448 N$24896 N$24895 "Straight Waveguide" sch_x=-173 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12449 N$24898 N$24897 "Straight Waveguide" sch_x=-173 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12450 N$24900 N$24899 "Straight Waveguide" sch_x=-173 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12451 N$24902 N$24901 "Straight Waveguide" sch_x=-173 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12452 N$24904 N$24903 "Straight Waveguide" sch_x=-173 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12453 N$24906 N$24905 "Straight Waveguide" sch_x=-173 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12454 N$24908 N$24907 "Straight Waveguide" sch_x=-173 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12455 N$24910 N$24909 "Straight Waveguide" sch_x=-173 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12456 N$24912 N$24911 "Straight Waveguide" sch_x=-173 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12457 N$24914 N$24913 "Straight Waveguide" sch_x=-173 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12458 N$24916 N$24915 "Straight Waveguide" sch_x=-173 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12459 N$24918 N$24917 "Straight Waveguide" sch_x=-173 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12460 N$24920 N$24919 "Straight Waveguide" sch_x=-173 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12461 N$24922 N$24921 "Straight Waveguide" sch_x=-173 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12462 N$24924 N$24923 "Straight Waveguide" sch_x=-173 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12463 N$24926 N$24925 "Straight Waveguide" sch_x=-173 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12464 N$24928 N$24927 "Straight Waveguide" sch_x=-173 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12465 N$24930 N$24929 "Straight Waveguide" sch_x=-173 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12466 N$24932 N$24931 "Straight Waveguide" sch_x=-173 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12467 N$24934 N$24933 "Straight Waveguide" sch_x=-173 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12468 N$24936 N$24935 "Straight Waveguide" sch_x=-173 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12469 N$24938 N$24937 "Straight Waveguide" sch_x=-173 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12470 N$24940 N$24939 "Straight Waveguide" sch_x=-173 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12471 N$24942 N$24941 "Straight Waveguide" sch_x=-173 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12472 N$24944 N$24943 "Straight Waveguide" sch_x=-173 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12473 N$24946 N$24945 "Straight Waveguide" sch_x=-173 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12474 N$24948 N$24947 "Straight Waveguide" sch_x=-173 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12475 N$24950 N$24949 "Straight Waveguide" sch_x=-173 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12476 N$24952 N$24951 "Straight Waveguide" sch_x=-173 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12477 N$24954 N$24953 "Straight Waveguide" sch_x=-173 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12478 N$24956 N$24955 "Straight Waveguide" sch_x=-173 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12479 N$24958 N$24957 "Straight Waveguide" sch_x=-173 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12480 N$24960 N$24959 "Straight Waveguide" sch_x=-173 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12481 N$24962 N$24961 "Straight Waveguide" sch_x=-173 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12482 N$24964 N$24963 "Straight Waveguide" sch_x=-173 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12483 N$24966 N$24965 "Straight Waveguide" sch_x=-173 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12484 N$24968 N$24967 "Straight Waveguide" sch_x=-173 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12485 N$24970 N$24969 "Straight Waveguide" sch_x=-173 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12486 N$24972 N$24971 "Straight Waveguide" sch_x=-173 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12487 N$24974 N$24973 "Straight Waveguide" sch_x=-171 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12488 N$24976 N$24975 "Straight Waveguide" sch_x=-171 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12489 N$24978 N$24977 "Straight Waveguide" sch_x=-171 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12490 N$24980 N$24979 "Straight Waveguide" sch_x=-171 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12491 N$24982 N$24981 "Straight Waveguide" sch_x=-171 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12492 N$24984 N$24983 "Straight Waveguide" sch_x=-171 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12493 N$24986 N$24985 "Straight Waveguide" sch_x=-171 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12494 N$24988 N$24987 "Straight Waveguide" sch_x=-171 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12495 N$24990 N$24989 "Straight Waveguide" sch_x=-171 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12496 N$24992 N$24991 "Straight Waveguide" sch_x=-171 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12497 N$24994 N$24993 "Straight Waveguide" sch_x=-171 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12498 N$24996 N$24995 "Straight Waveguide" sch_x=-171 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12499 N$24998 N$24997 "Straight Waveguide" sch_x=-171 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12500 N$25000 N$24999 "Straight Waveguide" sch_x=-171 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12501 N$25002 N$25001 "Straight Waveguide" sch_x=-171 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12502 N$25004 N$25003 "Straight Waveguide" sch_x=-171 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12503 N$25006 N$25005 "Straight Waveguide" sch_x=-171 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12504 N$25008 N$25007 "Straight Waveguide" sch_x=-171 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12505 N$25010 N$25009 "Straight Waveguide" sch_x=-171 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12506 N$25012 N$25011 "Straight Waveguide" sch_x=-171 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12507 N$25014 N$25013 "Straight Waveguide" sch_x=-171 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12508 N$25016 N$25015 "Straight Waveguide" sch_x=-171 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12509 N$25018 N$25017 "Straight Waveguide" sch_x=-171 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12510 N$25020 N$25019 "Straight Waveguide" sch_x=-171 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12511 N$25022 N$25021 "Straight Waveguide" sch_x=-171 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12512 N$25024 N$25023 "Straight Waveguide" sch_x=-171 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12513 N$25026 N$25025 "Straight Waveguide" sch_x=-171 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12514 N$25028 N$25027 "Straight Waveguide" sch_x=-171 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12515 N$25030 N$25029 "Straight Waveguide" sch_x=-171 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12516 N$25032 N$25031 "Straight Waveguide" sch_x=-171 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12517 N$25034 N$25033 "Straight Waveguide" sch_x=-171 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12518 N$25036 N$25035 "Straight Waveguide" sch_x=-171 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12519 N$25038 N$25037 "Straight Waveguide" sch_x=-171 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12520 N$25040 N$25039 "Straight Waveguide" sch_x=-171 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12521 N$25042 N$25041 "Straight Waveguide" sch_x=-171 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12522 N$25044 N$25043 "Straight Waveguide" sch_x=-171 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12523 N$25046 N$25045 "Straight Waveguide" sch_x=-171 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12524 N$25048 N$25047 "Straight Waveguide" sch_x=-171 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12525 N$25050 N$25049 "Straight Waveguide" sch_x=-171 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12526 N$25052 N$25051 "Straight Waveguide" sch_x=-171 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12527 N$25054 N$25053 "Straight Waveguide" sch_x=-171 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12528 N$25056 N$25055 "Straight Waveguide" sch_x=-171 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12529 N$25058 N$25057 "Straight Waveguide" sch_x=-171 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12530 N$25060 N$25059 "Straight Waveguide" sch_x=-171 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12531 N$25062 N$25061 "Straight Waveguide" sch_x=-169 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12532 N$25064 N$25063 "Straight Waveguide" sch_x=-169 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12533 N$25066 N$25065 "Straight Waveguide" sch_x=-169 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12534 N$25068 N$25067 "Straight Waveguide" sch_x=-169 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12535 N$25070 N$25069 "Straight Waveguide" sch_x=-169 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12536 N$25072 N$25071 "Straight Waveguide" sch_x=-169 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12537 N$25074 N$25073 "Straight Waveguide" sch_x=-169 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12538 N$25076 N$25075 "Straight Waveguide" sch_x=-169 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12539 N$25078 N$25077 "Straight Waveguide" sch_x=-169 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12540 N$25080 N$25079 "Straight Waveguide" sch_x=-169 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12541 N$25082 N$25081 "Straight Waveguide" sch_x=-169 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12542 N$25084 N$25083 "Straight Waveguide" sch_x=-169 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12543 N$25086 N$25085 "Straight Waveguide" sch_x=-169 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12544 N$25088 N$25087 "Straight Waveguide" sch_x=-169 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12545 N$25090 N$25089 "Straight Waveguide" sch_x=-169 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12546 N$25092 N$25091 "Straight Waveguide" sch_x=-169 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12547 N$25094 N$25093 "Straight Waveguide" sch_x=-169 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12548 N$25096 N$25095 "Straight Waveguide" sch_x=-169 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12549 N$25098 N$25097 "Straight Waveguide" sch_x=-169 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12550 N$25100 N$25099 "Straight Waveguide" sch_x=-169 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12551 N$25102 N$25101 "Straight Waveguide" sch_x=-169 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12552 N$25104 N$25103 "Straight Waveguide" sch_x=-169 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12553 N$25106 N$25105 "Straight Waveguide" sch_x=-169 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12554 N$25108 N$25107 "Straight Waveguide" sch_x=-169 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12555 N$25110 N$25109 "Straight Waveguide" sch_x=-169 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12556 N$25112 N$25111 "Straight Waveguide" sch_x=-169 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12557 N$25114 N$25113 "Straight Waveguide" sch_x=-169 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12558 N$25116 N$25115 "Straight Waveguide" sch_x=-169 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12559 N$25118 N$25117 "Straight Waveguide" sch_x=-169 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12560 N$25120 N$25119 "Straight Waveguide" sch_x=-169 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12561 N$25122 N$25121 "Straight Waveguide" sch_x=-169 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12562 N$25124 N$25123 "Straight Waveguide" sch_x=-169 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12563 N$25126 N$25125 "Straight Waveguide" sch_x=-169 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12564 N$25128 N$25127 "Straight Waveguide" sch_x=-169 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12565 N$25130 N$25129 "Straight Waveguide" sch_x=-169 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12566 N$25132 N$25131 "Straight Waveguide" sch_x=-169 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12567 N$25134 N$25133 "Straight Waveguide" sch_x=-169 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12568 N$25136 N$25135 "Straight Waveguide" sch_x=-169 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12569 N$25138 N$25137 "Straight Waveguide" sch_x=-169 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12570 N$25140 N$25139 "Straight Waveguide" sch_x=-169 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12571 N$25142 N$25141 "Straight Waveguide" sch_x=-169 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12572 N$25144 N$25143 "Straight Waveguide" sch_x=-169 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12573 N$25146 N$25145 "Straight Waveguide" sch_x=-167 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12574 N$25148 N$25147 "Straight Waveguide" sch_x=-167 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12575 N$25150 N$25149 "Straight Waveguide" sch_x=-167 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12576 N$25152 N$25151 "Straight Waveguide" sch_x=-167 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12577 N$25154 N$25153 "Straight Waveguide" sch_x=-167 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12578 N$25156 N$25155 "Straight Waveguide" sch_x=-167 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12579 N$25158 N$25157 "Straight Waveguide" sch_x=-167 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12580 N$25160 N$25159 "Straight Waveguide" sch_x=-167 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12581 N$25162 N$25161 "Straight Waveguide" sch_x=-167 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12582 N$25164 N$25163 "Straight Waveguide" sch_x=-167 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12583 N$25166 N$25165 "Straight Waveguide" sch_x=-167 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12584 N$25168 N$25167 "Straight Waveguide" sch_x=-167 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12585 N$25170 N$25169 "Straight Waveguide" sch_x=-167 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12586 N$25172 N$25171 "Straight Waveguide" sch_x=-167 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12587 N$25174 N$25173 "Straight Waveguide" sch_x=-167 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12588 N$25176 N$25175 "Straight Waveguide" sch_x=-167 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12589 N$25178 N$25177 "Straight Waveguide" sch_x=-167 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12590 N$25180 N$25179 "Straight Waveguide" sch_x=-167 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12591 N$25182 N$25181 "Straight Waveguide" sch_x=-167 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12592 N$25184 N$25183 "Straight Waveguide" sch_x=-167 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12593 N$25186 N$25185 "Straight Waveguide" sch_x=-167 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12594 N$25188 N$25187 "Straight Waveguide" sch_x=-167 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12595 N$25190 N$25189 "Straight Waveguide" sch_x=-167 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12596 N$25192 N$25191 "Straight Waveguide" sch_x=-167 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12597 N$25194 N$25193 "Straight Waveguide" sch_x=-167 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12598 N$25196 N$25195 "Straight Waveguide" sch_x=-167 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12599 N$25198 N$25197 "Straight Waveguide" sch_x=-167 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12600 N$25200 N$25199 "Straight Waveguide" sch_x=-167 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12601 N$25202 N$25201 "Straight Waveguide" sch_x=-167 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12602 N$25204 N$25203 "Straight Waveguide" sch_x=-167 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12603 N$25206 N$25205 "Straight Waveguide" sch_x=-167 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12604 N$25208 N$25207 "Straight Waveguide" sch_x=-167 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12605 N$25210 N$25209 "Straight Waveguide" sch_x=-167 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12606 N$25212 N$25211 "Straight Waveguide" sch_x=-167 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12607 N$25214 N$25213 "Straight Waveguide" sch_x=-167 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12608 N$25216 N$25215 "Straight Waveguide" sch_x=-167 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12609 N$25218 N$25217 "Straight Waveguide" sch_x=-167 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12610 N$25220 N$25219 "Straight Waveguide" sch_x=-167 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12611 N$25222 N$25221 "Straight Waveguide" sch_x=-167 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12612 N$25224 N$25223 "Straight Waveguide" sch_x=-167 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12613 N$25226 N$25225 "Straight Waveguide" sch_x=-165 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12614 N$25228 N$25227 "Straight Waveguide" sch_x=-165 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12615 N$25230 N$25229 "Straight Waveguide" sch_x=-165 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12616 N$25232 N$25231 "Straight Waveguide" sch_x=-165 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12617 N$25234 N$25233 "Straight Waveguide" sch_x=-165 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12618 N$25236 N$25235 "Straight Waveguide" sch_x=-165 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12619 N$25238 N$25237 "Straight Waveguide" sch_x=-165 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12620 N$25240 N$25239 "Straight Waveguide" sch_x=-165 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12621 N$25242 N$25241 "Straight Waveguide" sch_x=-165 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12622 N$25244 N$25243 "Straight Waveguide" sch_x=-165 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12623 N$25246 N$25245 "Straight Waveguide" sch_x=-165 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12624 N$25248 N$25247 "Straight Waveguide" sch_x=-165 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12625 N$25250 N$25249 "Straight Waveguide" sch_x=-165 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12626 N$25252 N$25251 "Straight Waveguide" sch_x=-165 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12627 N$25254 N$25253 "Straight Waveguide" sch_x=-165 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12628 N$25256 N$25255 "Straight Waveguide" sch_x=-165 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12629 N$25258 N$25257 "Straight Waveguide" sch_x=-165 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12630 N$25260 N$25259 "Straight Waveguide" sch_x=-165 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12631 N$25262 N$25261 "Straight Waveguide" sch_x=-165 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12632 N$25264 N$25263 "Straight Waveguide" sch_x=-165 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12633 N$25266 N$25265 "Straight Waveguide" sch_x=-165 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12634 N$25268 N$25267 "Straight Waveguide" sch_x=-165 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12635 N$25270 N$25269 "Straight Waveguide" sch_x=-165 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12636 N$25272 N$25271 "Straight Waveguide" sch_x=-165 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12637 N$25274 N$25273 "Straight Waveguide" sch_x=-165 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12638 N$25276 N$25275 "Straight Waveguide" sch_x=-165 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12639 N$25278 N$25277 "Straight Waveguide" sch_x=-165 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12640 N$25280 N$25279 "Straight Waveguide" sch_x=-165 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12641 N$25282 N$25281 "Straight Waveguide" sch_x=-165 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12642 N$25284 N$25283 "Straight Waveguide" sch_x=-165 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12643 N$25286 N$25285 "Straight Waveguide" sch_x=-165 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12644 N$25288 N$25287 "Straight Waveguide" sch_x=-165 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12645 N$25290 N$25289 "Straight Waveguide" sch_x=-165 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12646 N$25292 N$25291 "Straight Waveguide" sch_x=-165 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12647 N$25294 N$25293 "Straight Waveguide" sch_x=-165 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12648 N$25296 N$25295 "Straight Waveguide" sch_x=-165 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12649 N$25298 N$25297 "Straight Waveguide" sch_x=-165 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12650 N$25300 N$25299 "Straight Waveguide" sch_x=-165 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12651 N$25302 N$25301 "Straight Waveguide" sch_x=-163 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12652 N$25304 N$25303 "Straight Waveguide" sch_x=-163 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12653 N$25306 N$25305 "Straight Waveguide" sch_x=-163 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12654 N$25308 N$25307 "Straight Waveguide" sch_x=-163 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12655 N$25310 N$25309 "Straight Waveguide" sch_x=-163 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12656 N$25312 N$25311 "Straight Waveguide" sch_x=-163 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12657 N$25314 N$25313 "Straight Waveguide" sch_x=-163 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12658 N$25316 N$25315 "Straight Waveguide" sch_x=-163 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12659 N$25318 N$25317 "Straight Waveguide" sch_x=-163 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12660 N$25320 N$25319 "Straight Waveguide" sch_x=-163 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12661 N$25322 N$25321 "Straight Waveguide" sch_x=-163 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12662 N$25324 N$25323 "Straight Waveguide" sch_x=-163 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12663 N$25326 N$25325 "Straight Waveguide" sch_x=-163 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12664 N$25328 N$25327 "Straight Waveguide" sch_x=-163 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12665 N$25330 N$25329 "Straight Waveguide" sch_x=-163 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12666 N$25332 N$25331 "Straight Waveguide" sch_x=-163 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12667 N$25334 N$25333 "Straight Waveguide" sch_x=-163 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12668 N$25336 N$25335 "Straight Waveguide" sch_x=-163 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12669 N$25338 N$25337 "Straight Waveguide" sch_x=-163 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12670 N$25340 N$25339 "Straight Waveguide" sch_x=-163 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12671 N$25342 N$25341 "Straight Waveguide" sch_x=-163 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12672 N$25344 N$25343 "Straight Waveguide" sch_x=-163 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12673 N$25346 N$25345 "Straight Waveguide" sch_x=-163 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12674 N$25348 N$25347 "Straight Waveguide" sch_x=-163 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12675 N$25350 N$25349 "Straight Waveguide" sch_x=-163 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12676 N$25352 N$25351 "Straight Waveguide" sch_x=-163 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12677 N$25354 N$25353 "Straight Waveguide" sch_x=-163 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12678 N$25356 N$25355 "Straight Waveguide" sch_x=-163 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12679 N$25358 N$25357 "Straight Waveguide" sch_x=-163 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12680 N$25360 N$25359 "Straight Waveguide" sch_x=-163 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12681 N$25362 N$25361 "Straight Waveguide" sch_x=-163 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12682 N$25364 N$25363 "Straight Waveguide" sch_x=-163 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12683 N$25366 N$25365 "Straight Waveguide" sch_x=-163 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12684 N$25368 N$25367 "Straight Waveguide" sch_x=-163 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12685 N$25370 N$25369 "Straight Waveguide" sch_x=-163 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12686 N$25372 N$25371 "Straight Waveguide" sch_x=-163 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12687 N$25374 N$25373 "Straight Waveguide" sch_x=-161 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12688 N$25376 N$25375 "Straight Waveguide" sch_x=-161 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12689 N$25378 N$25377 "Straight Waveguide" sch_x=-161 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12690 N$25380 N$25379 "Straight Waveguide" sch_x=-161 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12691 N$25382 N$25381 "Straight Waveguide" sch_x=-161 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12692 N$25384 N$25383 "Straight Waveguide" sch_x=-161 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12693 N$25386 N$25385 "Straight Waveguide" sch_x=-161 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12694 N$25388 N$25387 "Straight Waveguide" sch_x=-161 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12695 N$25390 N$25389 "Straight Waveguide" sch_x=-161 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12696 N$25392 N$25391 "Straight Waveguide" sch_x=-161 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12697 N$25394 N$25393 "Straight Waveguide" sch_x=-161 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12698 N$25396 N$25395 "Straight Waveguide" sch_x=-161 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12699 N$25398 N$25397 "Straight Waveguide" sch_x=-161 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12700 N$25400 N$25399 "Straight Waveguide" sch_x=-161 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12701 N$25402 N$25401 "Straight Waveguide" sch_x=-161 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12702 N$25404 N$25403 "Straight Waveguide" sch_x=-161 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12703 N$25406 N$25405 "Straight Waveguide" sch_x=-161 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12704 N$25408 N$25407 "Straight Waveguide" sch_x=-161 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12705 N$25410 N$25409 "Straight Waveguide" sch_x=-161 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12706 N$25412 N$25411 "Straight Waveguide" sch_x=-161 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12707 N$25414 N$25413 "Straight Waveguide" sch_x=-161 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12708 N$25416 N$25415 "Straight Waveguide" sch_x=-161 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12709 N$25418 N$25417 "Straight Waveguide" sch_x=-161 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12710 N$25420 N$25419 "Straight Waveguide" sch_x=-161 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12711 N$25422 N$25421 "Straight Waveguide" sch_x=-161 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12712 N$25424 N$25423 "Straight Waveguide" sch_x=-161 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12713 N$25426 N$25425 "Straight Waveguide" sch_x=-161 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12714 N$25428 N$25427 "Straight Waveguide" sch_x=-161 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12715 N$25430 N$25429 "Straight Waveguide" sch_x=-161 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12716 N$25432 N$25431 "Straight Waveguide" sch_x=-161 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12717 N$25434 N$25433 "Straight Waveguide" sch_x=-161 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12718 N$25436 N$25435 "Straight Waveguide" sch_x=-161 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12719 N$25438 N$25437 "Straight Waveguide" sch_x=-161 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12720 N$25440 N$25439 "Straight Waveguide" sch_x=-161 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12721 N$25442 N$25441 "Straight Waveguide" sch_x=-159 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12722 N$25444 N$25443 "Straight Waveguide" sch_x=-159 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12723 N$25446 N$25445 "Straight Waveguide" sch_x=-159 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12724 N$25448 N$25447 "Straight Waveguide" sch_x=-159 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12725 N$25450 N$25449 "Straight Waveguide" sch_x=-159 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12726 N$25452 N$25451 "Straight Waveguide" sch_x=-159 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12727 N$25454 N$25453 "Straight Waveguide" sch_x=-159 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12728 N$25456 N$25455 "Straight Waveguide" sch_x=-159 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12729 N$25458 N$25457 "Straight Waveguide" sch_x=-159 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12730 N$25460 N$25459 "Straight Waveguide" sch_x=-159 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12731 N$25462 N$25461 "Straight Waveguide" sch_x=-159 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12732 N$25464 N$25463 "Straight Waveguide" sch_x=-159 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12733 N$25466 N$25465 "Straight Waveguide" sch_x=-159 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12734 N$25468 N$25467 "Straight Waveguide" sch_x=-159 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12735 N$25470 N$25469 "Straight Waveguide" sch_x=-159 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12736 N$25472 N$25471 "Straight Waveguide" sch_x=-159 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12737 N$25474 N$25473 "Straight Waveguide" sch_x=-159 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12738 N$25476 N$25475 "Straight Waveguide" sch_x=-159 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12739 N$25478 N$25477 "Straight Waveguide" sch_x=-159 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12740 N$25480 N$25479 "Straight Waveguide" sch_x=-159 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12741 N$25482 N$25481 "Straight Waveguide" sch_x=-159 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12742 N$25484 N$25483 "Straight Waveguide" sch_x=-159 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12743 N$25486 N$25485 "Straight Waveguide" sch_x=-159 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12744 N$25488 N$25487 "Straight Waveguide" sch_x=-159 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12745 N$25490 N$25489 "Straight Waveguide" sch_x=-159 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12746 N$25492 N$25491 "Straight Waveguide" sch_x=-159 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12747 N$25494 N$25493 "Straight Waveguide" sch_x=-159 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12748 N$25496 N$25495 "Straight Waveguide" sch_x=-159 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12749 N$25498 N$25497 "Straight Waveguide" sch_x=-159 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12750 N$25500 N$25499 "Straight Waveguide" sch_x=-159 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12751 N$25502 N$25501 "Straight Waveguide" sch_x=-159 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12752 N$25504 N$25503 "Straight Waveguide" sch_x=-159 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12753 N$25506 N$25505 "Straight Waveguide" sch_x=-157 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12754 N$25508 N$25507 "Straight Waveguide" sch_x=-157 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12755 N$25510 N$25509 "Straight Waveguide" sch_x=-157 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12756 N$25512 N$25511 "Straight Waveguide" sch_x=-157 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12757 N$25514 N$25513 "Straight Waveguide" sch_x=-157 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12758 N$25516 N$25515 "Straight Waveguide" sch_x=-157 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12759 N$25518 N$25517 "Straight Waveguide" sch_x=-157 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12760 N$25520 N$25519 "Straight Waveguide" sch_x=-157 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12761 N$25522 N$25521 "Straight Waveguide" sch_x=-157 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12762 N$25524 N$25523 "Straight Waveguide" sch_x=-157 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12763 N$25526 N$25525 "Straight Waveguide" sch_x=-157 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12764 N$25528 N$25527 "Straight Waveguide" sch_x=-157 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12765 N$25530 N$25529 "Straight Waveguide" sch_x=-157 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12766 N$25532 N$25531 "Straight Waveguide" sch_x=-157 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12767 N$25534 N$25533 "Straight Waveguide" sch_x=-157 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12768 N$25536 N$25535 "Straight Waveguide" sch_x=-157 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12769 N$25538 N$25537 "Straight Waveguide" sch_x=-157 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12770 N$25540 N$25539 "Straight Waveguide" sch_x=-157 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12771 N$25542 N$25541 "Straight Waveguide" sch_x=-157 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12772 N$25544 N$25543 "Straight Waveguide" sch_x=-157 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12773 N$25546 N$25545 "Straight Waveguide" sch_x=-157 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12774 N$25548 N$25547 "Straight Waveguide" sch_x=-157 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12775 N$25550 N$25549 "Straight Waveguide" sch_x=-157 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12776 N$25552 N$25551 "Straight Waveguide" sch_x=-157 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12777 N$25554 N$25553 "Straight Waveguide" sch_x=-157 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12778 N$25556 N$25555 "Straight Waveguide" sch_x=-157 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12779 N$25558 N$25557 "Straight Waveguide" sch_x=-157 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12780 N$25560 N$25559 "Straight Waveguide" sch_x=-157 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12781 N$25562 N$25561 "Straight Waveguide" sch_x=-157 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12782 N$25564 N$25563 "Straight Waveguide" sch_x=-157 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12783 N$25566 N$25565 "Straight Waveguide" sch_x=-155 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12784 N$25568 N$25567 "Straight Waveguide" sch_x=-155 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12785 N$25570 N$25569 "Straight Waveguide" sch_x=-155 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12786 N$25572 N$25571 "Straight Waveguide" sch_x=-155 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12787 N$25574 N$25573 "Straight Waveguide" sch_x=-155 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12788 N$25576 N$25575 "Straight Waveguide" sch_x=-155 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12789 N$25578 N$25577 "Straight Waveguide" sch_x=-155 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12790 N$25580 N$25579 "Straight Waveguide" sch_x=-155 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12791 N$25582 N$25581 "Straight Waveguide" sch_x=-155 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12792 N$25584 N$25583 "Straight Waveguide" sch_x=-155 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12793 N$25586 N$25585 "Straight Waveguide" sch_x=-155 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12794 N$25588 N$25587 "Straight Waveguide" sch_x=-155 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12795 N$25590 N$25589 "Straight Waveguide" sch_x=-155 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12796 N$25592 N$25591 "Straight Waveguide" sch_x=-155 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12797 N$25594 N$25593 "Straight Waveguide" sch_x=-155 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12798 N$25596 N$25595 "Straight Waveguide" sch_x=-155 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12799 N$25598 N$25597 "Straight Waveguide" sch_x=-155 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12800 N$25600 N$25599 "Straight Waveguide" sch_x=-155 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12801 N$25602 N$25601 "Straight Waveguide" sch_x=-155 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12802 N$25604 N$25603 "Straight Waveguide" sch_x=-155 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12803 N$25606 N$25605 "Straight Waveguide" sch_x=-155 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12804 N$25608 N$25607 "Straight Waveguide" sch_x=-155 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12805 N$25610 N$25609 "Straight Waveguide" sch_x=-155 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12806 N$25612 N$25611 "Straight Waveguide" sch_x=-155 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12807 N$25614 N$25613 "Straight Waveguide" sch_x=-155 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12808 N$25616 N$25615 "Straight Waveguide" sch_x=-155 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12809 N$25618 N$25617 "Straight Waveguide" sch_x=-155 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12810 N$25620 N$25619 "Straight Waveguide" sch_x=-155 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12811 N$25622 N$25621 "Straight Waveguide" sch_x=-153 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12812 N$25624 N$25623 "Straight Waveguide" sch_x=-153 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12813 N$25626 N$25625 "Straight Waveguide" sch_x=-153 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12814 N$25628 N$25627 "Straight Waveguide" sch_x=-153 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12815 N$25630 N$25629 "Straight Waveguide" sch_x=-153 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12816 N$25632 N$25631 "Straight Waveguide" sch_x=-153 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12817 N$25634 N$25633 "Straight Waveguide" sch_x=-153 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12818 N$25636 N$25635 "Straight Waveguide" sch_x=-153 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12819 N$25638 N$25637 "Straight Waveguide" sch_x=-153 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12820 N$25640 N$25639 "Straight Waveguide" sch_x=-153 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12821 N$25642 N$25641 "Straight Waveguide" sch_x=-153 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12822 N$25644 N$25643 "Straight Waveguide" sch_x=-153 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12823 N$25646 N$25645 "Straight Waveguide" sch_x=-153 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12824 N$25648 N$25647 "Straight Waveguide" sch_x=-153 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12825 N$25650 N$25649 "Straight Waveguide" sch_x=-153 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12826 N$25652 N$25651 "Straight Waveguide" sch_x=-153 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12827 N$25654 N$25653 "Straight Waveguide" sch_x=-153 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12828 N$25656 N$25655 "Straight Waveguide" sch_x=-153 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12829 N$25658 N$25657 "Straight Waveguide" sch_x=-153 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12830 N$25660 N$25659 "Straight Waveguide" sch_x=-153 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12831 N$25662 N$25661 "Straight Waveguide" sch_x=-153 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12832 N$25664 N$25663 "Straight Waveguide" sch_x=-153 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12833 N$25666 N$25665 "Straight Waveguide" sch_x=-153 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12834 N$25668 N$25667 "Straight Waveguide" sch_x=-153 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12835 N$25670 N$25669 "Straight Waveguide" sch_x=-153 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12836 N$25672 N$25671 "Straight Waveguide" sch_x=-153 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12837 N$25674 N$25673 "Straight Waveguide" sch_x=-151 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12838 N$25676 N$25675 "Straight Waveguide" sch_x=-151 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12839 N$25678 N$25677 "Straight Waveguide" sch_x=-151 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12840 N$25680 N$25679 "Straight Waveguide" sch_x=-151 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12841 N$25682 N$25681 "Straight Waveguide" sch_x=-151 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12842 N$25684 N$25683 "Straight Waveguide" sch_x=-151 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12843 N$25686 N$25685 "Straight Waveguide" sch_x=-151 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12844 N$25688 N$25687 "Straight Waveguide" sch_x=-151 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12845 N$25690 N$25689 "Straight Waveguide" sch_x=-151 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12846 N$25692 N$25691 "Straight Waveguide" sch_x=-151 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12847 N$25694 N$25693 "Straight Waveguide" sch_x=-151 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12848 N$25696 N$25695 "Straight Waveguide" sch_x=-151 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12849 N$25698 N$25697 "Straight Waveguide" sch_x=-151 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12850 N$25700 N$25699 "Straight Waveguide" sch_x=-151 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12851 N$25702 N$25701 "Straight Waveguide" sch_x=-151 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12852 N$25704 N$25703 "Straight Waveguide" sch_x=-151 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12853 N$25706 N$25705 "Straight Waveguide" sch_x=-151 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12854 N$25708 N$25707 "Straight Waveguide" sch_x=-151 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12855 N$25710 N$25709 "Straight Waveguide" sch_x=-151 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12856 N$25712 N$25711 "Straight Waveguide" sch_x=-151 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12857 N$25714 N$25713 "Straight Waveguide" sch_x=-151 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12858 N$25716 N$25715 "Straight Waveguide" sch_x=-151 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12859 N$25718 N$25717 "Straight Waveguide" sch_x=-151 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12860 N$25720 N$25719 "Straight Waveguide" sch_x=-151 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12861 N$25722 N$25721 "Straight Waveguide" sch_x=-149 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12862 N$25724 N$25723 "Straight Waveguide" sch_x=-149 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12863 N$25726 N$25725 "Straight Waveguide" sch_x=-149 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12864 N$25728 N$25727 "Straight Waveguide" sch_x=-149 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12865 N$25730 N$25729 "Straight Waveguide" sch_x=-149 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12866 N$25732 N$25731 "Straight Waveguide" sch_x=-149 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12867 N$25734 N$25733 "Straight Waveguide" sch_x=-149 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12868 N$25736 N$25735 "Straight Waveguide" sch_x=-149 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12869 N$25738 N$25737 "Straight Waveguide" sch_x=-149 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12870 N$25740 N$25739 "Straight Waveguide" sch_x=-149 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12871 N$25742 N$25741 "Straight Waveguide" sch_x=-149 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12872 N$25744 N$25743 "Straight Waveguide" sch_x=-149 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12873 N$25746 N$25745 "Straight Waveguide" sch_x=-149 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12874 N$25748 N$25747 "Straight Waveguide" sch_x=-149 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12875 N$25750 N$25749 "Straight Waveguide" sch_x=-149 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12876 N$25752 N$25751 "Straight Waveguide" sch_x=-149 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12877 N$25754 N$25753 "Straight Waveguide" sch_x=-149 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12878 N$25756 N$25755 "Straight Waveguide" sch_x=-149 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12879 N$25758 N$25757 "Straight Waveguide" sch_x=-149 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12880 N$25760 N$25759 "Straight Waveguide" sch_x=-149 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12881 N$25762 N$25761 "Straight Waveguide" sch_x=-149 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12882 N$25764 N$25763 "Straight Waveguide" sch_x=-149 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12883 N$25766 N$25765 "Straight Waveguide" sch_x=-147 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12884 N$25768 N$25767 "Straight Waveguide" sch_x=-147 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12885 N$25770 N$25769 "Straight Waveguide" sch_x=-147 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12886 N$25772 N$25771 "Straight Waveguide" sch_x=-147 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12887 N$25774 N$25773 "Straight Waveguide" sch_x=-147 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12888 N$25776 N$25775 "Straight Waveguide" sch_x=-147 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12889 N$25778 N$25777 "Straight Waveguide" sch_x=-147 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12890 N$25780 N$25779 "Straight Waveguide" sch_x=-147 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12891 N$25782 N$25781 "Straight Waveguide" sch_x=-147 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12892 N$25784 N$25783 "Straight Waveguide" sch_x=-147 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12893 N$25786 N$25785 "Straight Waveguide" sch_x=-147 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12894 N$25788 N$25787 "Straight Waveguide" sch_x=-147 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12895 N$25790 N$25789 "Straight Waveguide" sch_x=-147 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12896 N$25792 N$25791 "Straight Waveguide" sch_x=-147 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12897 N$25794 N$25793 "Straight Waveguide" sch_x=-147 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12898 N$25796 N$25795 "Straight Waveguide" sch_x=-147 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12899 N$25798 N$25797 "Straight Waveguide" sch_x=-147 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12900 N$25800 N$25799 "Straight Waveguide" sch_x=-147 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12901 N$25802 N$25801 "Straight Waveguide" sch_x=-147 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12902 N$25804 N$25803 "Straight Waveguide" sch_x=-147 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12903 N$25806 N$25805 "Straight Waveguide" sch_x=-145 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12904 N$25808 N$25807 "Straight Waveguide" sch_x=-145 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12905 N$25810 N$25809 "Straight Waveguide" sch_x=-145 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12906 N$25812 N$25811 "Straight Waveguide" sch_x=-145 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12907 N$25814 N$25813 "Straight Waveguide" sch_x=-145 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12908 N$25816 N$25815 "Straight Waveguide" sch_x=-145 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12909 N$25818 N$25817 "Straight Waveguide" sch_x=-145 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12910 N$25820 N$25819 "Straight Waveguide" sch_x=-145 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12911 N$25822 N$25821 "Straight Waveguide" sch_x=-145 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12912 N$25824 N$25823 "Straight Waveguide" sch_x=-145 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12913 N$25826 N$25825 "Straight Waveguide" sch_x=-145 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12914 N$25828 N$25827 "Straight Waveguide" sch_x=-145 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12915 N$25830 N$25829 "Straight Waveguide" sch_x=-145 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12916 N$25832 N$25831 "Straight Waveguide" sch_x=-145 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12917 N$25834 N$25833 "Straight Waveguide" sch_x=-145 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12918 N$25836 N$25835 "Straight Waveguide" sch_x=-145 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12919 N$25838 N$25837 "Straight Waveguide" sch_x=-145 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12920 N$25840 N$25839 "Straight Waveguide" sch_x=-145 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12921 N$25842 N$25841 "Straight Waveguide" sch_x=-143 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12922 N$25844 N$25843 "Straight Waveguide" sch_x=-143 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12923 N$25846 N$25845 "Straight Waveguide" sch_x=-143 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12924 N$25848 N$25847 "Straight Waveguide" sch_x=-143 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12925 N$25850 N$25849 "Straight Waveguide" sch_x=-143 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12926 N$25852 N$25851 "Straight Waveguide" sch_x=-143 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12927 N$25854 N$25853 "Straight Waveguide" sch_x=-143 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12928 N$25856 N$25855 "Straight Waveguide" sch_x=-143 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12929 N$25858 N$25857 "Straight Waveguide" sch_x=-143 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12930 N$25860 N$25859 "Straight Waveguide" sch_x=-143 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12931 N$25862 N$25861 "Straight Waveguide" sch_x=-143 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12932 N$25864 N$25863 "Straight Waveguide" sch_x=-143 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12933 N$25866 N$25865 "Straight Waveguide" sch_x=-143 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12934 N$25868 N$25867 "Straight Waveguide" sch_x=-143 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12935 N$25870 N$25869 "Straight Waveguide" sch_x=-143 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12936 N$25872 N$25871 "Straight Waveguide" sch_x=-143 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12937 N$25874 N$25873 "Straight Waveguide" sch_x=-141 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12938 N$25876 N$25875 "Straight Waveguide" sch_x=-141 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12939 N$25878 N$25877 "Straight Waveguide" sch_x=-141 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12940 N$25880 N$25879 "Straight Waveguide" sch_x=-141 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12941 N$25882 N$25881 "Straight Waveguide" sch_x=-141 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12942 N$25884 N$25883 "Straight Waveguide" sch_x=-141 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12943 N$25886 N$25885 "Straight Waveguide" sch_x=-141 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12944 N$25888 N$25887 "Straight Waveguide" sch_x=-141 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12945 N$25890 N$25889 "Straight Waveguide" sch_x=-141 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12946 N$25892 N$25891 "Straight Waveguide" sch_x=-141 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12947 N$25894 N$25893 "Straight Waveguide" sch_x=-141 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12948 N$25896 N$25895 "Straight Waveguide" sch_x=-141 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12949 N$25898 N$25897 "Straight Waveguide" sch_x=-141 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12950 N$25900 N$25899 "Straight Waveguide" sch_x=-141 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12951 N$25902 N$25901 "Straight Waveguide" sch_x=-139 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12952 N$25904 N$25903 "Straight Waveguide" sch_x=-139 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12953 N$25906 N$25905 "Straight Waveguide" sch_x=-139 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12954 N$25908 N$25907 "Straight Waveguide" sch_x=-139 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12955 N$25910 N$25909 "Straight Waveguide" sch_x=-139 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12956 N$25912 N$25911 "Straight Waveguide" sch_x=-139 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12957 N$25914 N$25913 "Straight Waveguide" sch_x=-139 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12958 N$25916 N$25915 "Straight Waveguide" sch_x=-139 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12959 N$25918 N$25917 "Straight Waveguide" sch_x=-139 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12960 N$25920 N$25919 "Straight Waveguide" sch_x=-139 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12961 N$25922 N$25921 "Straight Waveguide" sch_x=-139 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12962 N$25924 N$25923 "Straight Waveguide" sch_x=-139 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12963 N$25926 N$25925 "Straight Waveguide" sch_x=-137 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12964 N$25928 N$25927 "Straight Waveguide" sch_x=-137 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12965 N$25930 N$25929 "Straight Waveguide" sch_x=-137 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12966 N$25932 N$25931 "Straight Waveguide" sch_x=-137 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12967 N$25934 N$25933 "Straight Waveguide" sch_x=-137 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12968 N$25936 N$25935 "Straight Waveguide" sch_x=-137 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12969 N$25938 N$25937 "Straight Waveguide" sch_x=-137 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12970 N$25940 N$25939 "Straight Waveguide" sch_x=-137 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12971 N$25942 N$25941 "Straight Waveguide" sch_x=-137 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12972 N$25944 N$25943 "Straight Waveguide" sch_x=-137 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12973 N$25946 N$25945 "Straight Waveguide" sch_x=-135 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12974 N$25948 N$25947 "Straight Waveguide" sch_x=-135 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12975 N$25950 N$25949 "Straight Waveguide" sch_x=-135 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12976 N$25952 N$25951 "Straight Waveguide" sch_x=-135 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12977 N$25954 N$25953 "Straight Waveguide" sch_x=-135 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12978 N$25956 N$25955 "Straight Waveguide" sch_x=-135 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12979 N$25958 N$25957 "Straight Waveguide" sch_x=-135 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12980 N$25960 N$25959 "Straight Waveguide" sch_x=-135 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12981 N$25962 N$25961 "Straight Waveguide" sch_x=-133 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12982 N$25964 N$25963 "Straight Waveguide" sch_x=-133 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12983 N$25966 N$25965 "Straight Waveguide" sch_x=-133 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12984 N$25968 N$25967 "Straight Waveguide" sch_x=-133 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12985 N$25970 N$25969 "Straight Waveguide" sch_x=-133 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12986 N$25972 N$25971 "Straight Waveguide" sch_x=-133 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12987 N$25974 N$25973 "Straight Waveguide" sch_x=-131 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12988 N$25976 N$25975 "Straight Waveguide" sch_x=-131 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12989 N$25978 N$25977 "Straight Waveguide" sch_x=-131 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12990 N$25980 N$25979 "Straight Waveguide" sch_x=-131 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12991 N$25982 N$25981 "Straight Waveguide" sch_x=-129 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12992 N$25984 N$25983 "Straight Waveguide" sch_x=-129 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12993 N$25985 N$25986 "Straight Waveguide" sch_x=-189 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12994 N$25987 N$25988 "Straight Waveguide" sch_x=-188 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12995 N$25989 N$25990 "Straight Waveguide" sch_x=-187 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12996 N$25991 N$25992 "Straight Waveguide" sch_x=-186 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12997 N$25993 N$25994 "Straight Waveguide" sch_x=-185 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12998 N$25995 N$25996 "Straight Waveguide" sch_x=-184 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12999 N$25997 N$25998 "Straight Waveguide" sch_x=-183 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13000 N$25999 N$26000 "Straight Waveguide" sch_x=-182 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13001 N$26001 N$26002 "Straight Waveguide" sch_x=-181 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13002 N$26003 N$26004 "Straight Waveguide" sch_x=-180 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13003 N$26005 N$26006 "Straight Waveguide" sch_x=-179 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13004 N$26007 N$26008 "Straight Waveguide" sch_x=-178 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13005 N$26009 N$26010 "Straight Waveguide" sch_x=-177 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13006 N$26011 N$26012 "Straight Waveguide" sch_x=-176 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13007 N$26013 N$26014 "Straight Waveguide" sch_x=-175 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13008 N$26015 N$26016 "Straight Waveguide" sch_x=-174 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13009 N$26017 N$26018 "Straight Waveguide" sch_x=-173 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13010 N$26019 N$26020 "Straight Waveguide" sch_x=-172 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13011 N$26021 N$26022 "Straight Waveguide" sch_x=-171 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13012 N$26023 N$26024 "Straight Waveguide" sch_x=-170 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13013 N$26025 N$26026 "Straight Waveguide" sch_x=-169 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13014 N$26027 N$26028 "Straight Waveguide" sch_x=-168 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13015 N$26029 N$26030 "Straight Waveguide" sch_x=-167 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13016 N$26031 N$26032 "Straight Waveguide" sch_x=-166 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13017 N$26033 N$26034 "Straight Waveguide" sch_x=-165 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13018 N$26035 N$26036 "Straight Waveguide" sch_x=-164 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13019 N$26037 N$26038 "Straight Waveguide" sch_x=-163 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13020 N$26039 N$26040 "Straight Waveguide" sch_x=-162 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13021 N$26041 N$26042 "Straight Waveguide" sch_x=-161 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13022 N$26043 N$26044 "Straight Waveguide" sch_x=-160 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13023 N$26045 N$26046 "Straight Waveguide" sch_x=-159 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13024 N$26047 N$26048 "Straight Waveguide" sch_x=-158 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13025 N$26049 N$26050 "Straight Waveguide" sch_x=-157 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13026 N$26051 N$26052 "Straight Waveguide" sch_x=-156 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13027 N$26053 N$26054 "Straight Waveguide" sch_x=-155 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13028 N$26055 N$26056 "Straight Waveguide" sch_x=-154 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13029 N$26057 N$26058 "Straight Waveguide" sch_x=-153 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13030 N$26059 N$26060 "Straight Waveguide" sch_x=-152 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13031 N$26061 N$26062 "Straight Waveguide" sch_x=-151 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13032 N$26063 N$26064 "Straight Waveguide" sch_x=-150 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13033 N$26065 N$26066 "Straight Waveguide" sch_x=-149 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13034 N$26067 N$26068 "Straight Waveguide" sch_x=-148 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13035 N$26069 N$26070 "Straight Waveguide" sch_x=-147 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13036 N$26071 N$26072 "Straight Waveguide" sch_x=-146 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13037 N$26073 N$26074 "Straight Waveguide" sch_x=-145 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13038 N$26075 N$26076 "Straight Waveguide" sch_x=-144 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13039 N$26077 N$26078 "Straight Waveguide" sch_x=-143 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13040 N$26079 N$26080 "Straight Waveguide" sch_x=-142 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13041 N$26081 N$26082 "Straight Waveguide" sch_x=-141 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13042 N$26083 N$26084 "Straight Waveguide" sch_x=-140 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13043 N$26085 N$26086 "Straight Waveguide" sch_x=-139 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13044 N$26087 N$26088 "Straight Waveguide" sch_x=-138 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13045 N$26089 N$26090 "Straight Waveguide" sch_x=-137 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13046 N$26091 N$26092 "Straight Waveguide" sch_x=-136 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13047 N$26093 N$26094 "Straight Waveguide" sch_x=-135 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13048 N$26095 N$26096 "Straight Waveguide" sch_x=-134 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13049 N$26097 N$26098 "Straight Waveguide" sch_x=-133 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13050 N$26099 N$26100 "Straight Waveguide" sch_x=-132 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13051 N$26101 N$26102 "Straight Waveguide" sch_x=-131 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13052 N$26103 N$26104 "Straight Waveguide" sch_x=-130 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13053 N$26105 N$26106 "Straight Waveguide" sch_x=-129 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13054 N$26107 N$26108 "Straight Waveguide" sch_x=-128 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13055 N$26109 N$26110 "Straight Waveguide" sch_x=-127 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13056 N$26111 N$26112 "Straight Waveguide" sch_x=-127 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13057 N$26113 N$26114 "Straight Waveguide" sch_x=-128 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13058 N$26115 N$26116 "Straight Waveguide" sch_x=-129 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13059 N$26117 N$26118 "Straight Waveguide" sch_x=-130 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13060 N$26119 N$26120 "Straight Waveguide" sch_x=-131 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13061 N$26121 N$26122 "Straight Waveguide" sch_x=-132 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13062 N$26123 N$26124 "Straight Waveguide" sch_x=-133 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13063 N$26125 N$26126 "Straight Waveguide" sch_x=-134 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13064 N$26127 N$26128 "Straight Waveguide" sch_x=-135 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13065 N$26129 N$26130 "Straight Waveguide" sch_x=-136 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13066 N$26131 N$26132 "Straight Waveguide" sch_x=-137 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13067 N$26133 N$26134 "Straight Waveguide" sch_x=-138 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13068 N$26135 N$26136 "Straight Waveguide" sch_x=-139 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13069 N$26137 N$26138 "Straight Waveguide" sch_x=-140 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13070 N$26139 N$26140 "Straight Waveguide" sch_x=-141 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13071 N$26141 N$26142 "Straight Waveguide" sch_x=-142 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13072 N$26143 N$26144 "Straight Waveguide" sch_x=-143 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13073 N$26145 N$26146 "Straight Waveguide" sch_x=-144 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13074 N$26147 N$26148 "Straight Waveguide" sch_x=-145 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13075 N$26149 N$26150 "Straight Waveguide" sch_x=-146 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13076 N$26151 N$26152 "Straight Waveguide" sch_x=-147 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13077 N$26153 N$26154 "Straight Waveguide" sch_x=-148 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13078 N$26155 N$26156 "Straight Waveguide" sch_x=-149 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13079 N$26157 N$26158 "Straight Waveguide" sch_x=-150 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13080 N$26159 N$26160 "Straight Waveguide" sch_x=-151 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13081 N$26161 N$26162 "Straight Waveguide" sch_x=-152 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13082 N$26163 N$26164 "Straight Waveguide" sch_x=-153 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13083 N$26165 N$26166 "Straight Waveguide" sch_x=-154 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13084 N$26167 N$26168 "Straight Waveguide" sch_x=-155 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13085 N$26169 N$26170 "Straight Waveguide" sch_x=-156 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13086 N$26171 N$26172 "Straight Waveguide" sch_x=-157 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13087 N$26173 N$26174 "Straight Waveguide" sch_x=-158 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13088 N$26175 N$26176 "Straight Waveguide" sch_x=-159 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13089 N$26177 N$26178 "Straight Waveguide" sch_x=-160 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13090 N$26179 N$26180 "Straight Waveguide" sch_x=-161 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13091 N$26181 N$26182 "Straight Waveguide" sch_x=-162 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13092 N$26183 N$26184 "Straight Waveguide" sch_x=-163 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13093 N$26185 N$26186 "Straight Waveguide" sch_x=-164 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13094 N$26187 N$26188 "Straight Waveguide" sch_x=-165 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13095 N$26189 N$26190 "Straight Waveguide" sch_x=-166 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13096 N$26191 N$26192 "Straight Waveguide" sch_x=-167 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13097 N$26193 N$26194 "Straight Waveguide" sch_x=-168 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13098 N$26195 N$26196 "Straight Waveguide" sch_x=-169 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13099 N$26197 N$26198 "Straight Waveguide" sch_x=-170 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13100 N$26199 N$26200 "Straight Waveguide" sch_x=-171 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13101 N$26201 N$26202 "Straight Waveguide" sch_x=-172 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13102 N$26203 N$26204 "Straight Waveguide" sch_x=-173 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13103 N$26205 N$26206 "Straight Waveguide" sch_x=-174 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13104 N$26207 N$26208 "Straight Waveguide" sch_x=-175 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13105 N$26209 N$26210 "Straight Waveguide" sch_x=-176 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13106 N$26211 N$26212 "Straight Waveguide" sch_x=-177 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13107 N$26213 N$26214 "Straight Waveguide" sch_x=-178 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13108 N$26215 N$26216 "Straight Waveguide" sch_x=-179 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13109 N$26217 N$26218 "Straight Waveguide" sch_x=-180 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13110 N$26219 N$26220 "Straight Waveguide" sch_x=-181 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13111 N$26221 N$26222 "Straight Waveguide" sch_x=-182 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13112 N$26223 N$26224 "Straight Waveguide" sch_x=-183 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13113 N$26225 N$26226 "Straight Waveguide" sch_x=-184 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13114 N$26227 N$26228 "Straight Waveguide" sch_x=-185 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13115 N$26229 N$26230 "Straight Waveguide" sch_x=-186 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13116 N$26231 N$26232 "Straight Waveguide" sch_x=-187 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13117 N$26233 N$26234 "Straight Waveguide" sch_x=-188 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13118 N$26235 N$26236 "Straight Waveguide" sch_x=-189 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13119 N$26237 N$26238 "Straight Waveguide" sch_x=-190 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13120 N$26239 N$26240 "Straight Waveguide" sch_x=-190 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13121 N$26241 N$26242 "Straight Waveguide" sch_x=253 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13122 N$26243 N$26244 "Straight Waveguide" sch_x=253 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13123 N$26245 N$26246 "Straight Waveguide" sch_x=253 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13124 N$26247 N$26248 "Straight Waveguide" sch_x=253 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13125 N$26249 N$26250 "Straight Waveguide" sch_x=253 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13126 N$26251 N$26252 "Straight Waveguide" sch_x=253 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13127 N$26253 N$26254 "Straight Waveguide" sch_x=253 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13128 N$26255 N$26256 "Straight Waveguide" sch_x=253 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13129 N$26257 N$26258 "Straight Waveguide" sch_x=253 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13130 N$26259 N$26260 "Straight Waveguide" sch_x=253 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13131 N$26261 N$26262 "Straight Waveguide" sch_x=253 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13132 N$26263 N$26264 "Straight Waveguide" sch_x=253 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13133 N$26265 N$26266 "Straight Waveguide" sch_x=253 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13134 N$26267 N$26268 "Straight Waveguide" sch_x=253 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13135 N$26269 N$26270 "Straight Waveguide" sch_x=253 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13136 N$26271 N$26272 "Straight Waveguide" sch_x=253 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13137 N$26273 N$26274 "Straight Waveguide" sch_x=253 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13138 N$26275 N$26276 "Straight Waveguide" sch_x=253 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13139 N$26277 N$26278 "Straight Waveguide" sch_x=253 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13140 N$26279 N$26280 "Straight Waveguide" sch_x=253 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13141 N$26281 N$26282 "Straight Waveguide" sch_x=253 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13142 N$26283 N$26284 "Straight Waveguide" sch_x=253 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13143 N$26285 N$26286 "Straight Waveguide" sch_x=253 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13144 N$26287 N$26288 "Straight Waveguide" sch_x=253 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13145 N$26289 N$26290 "Straight Waveguide" sch_x=253 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13146 N$26291 N$26292 "Straight Waveguide" sch_x=253 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13147 N$26293 N$26294 "Straight Waveguide" sch_x=253 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13148 N$26295 N$26296 "Straight Waveguide" sch_x=253 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13149 N$26297 N$26298 "Straight Waveguide" sch_x=253 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13150 N$26299 N$26300 "Straight Waveguide" sch_x=253 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13151 N$26301 N$26302 "Straight Waveguide" sch_x=253 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13152 N$26303 N$26304 "Straight Waveguide" sch_x=253 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13153 N$26305 N$26306 "Straight Waveguide" sch_x=253 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13154 N$26307 N$26308 "Straight Waveguide" sch_x=253 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13155 N$26309 N$26310 "Straight Waveguide" sch_x=253 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13156 N$26311 N$26312 "Straight Waveguide" sch_x=253 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13157 N$26313 N$26314 "Straight Waveguide" sch_x=253 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13158 N$26315 N$26316 "Straight Waveguide" sch_x=253 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13159 N$26317 N$26318 "Straight Waveguide" sch_x=253 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13160 N$26319 N$26320 "Straight Waveguide" sch_x=253 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13161 N$26321 N$26322 "Straight Waveguide" sch_x=253 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13162 N$26323 N$26324 "Straight Waveguide" sch_x=253 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13163 N$26325 N$26326 "Straight Waveguide" sch_x=253 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13164 N$26327 N$26328 "Straight Waveguide" sch_x=253 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13165 N$26329 N$26330 "Straight Waveguide" sch_x=253 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13166 N$26331 N$26332 "Straight Waveguide" sch_x=253 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13167 N$26333 N$26334 "Straight Waveguide" sch_x=253 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13168 N$26335 N$26336 "Straight Waveguide" sch_x=253 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13169 N$26337 N$26338 "Straight Waveguide" sch_x=253 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13170 N$26339 N$26340 "Straight Waveguide" sch_x=253 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13171 N$26341 N$26342 "Straight Waveguide" sch_x=253 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13172 N$26343 N$26344 "Straight Waveguide" sch_x=253 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13173 N$26345 N$26346 "Straight Waveguide" sch_x=253 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13174 N$26347 N$26348 "Straight Waveguide" sch_x=253 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13175 N$26349 N$26350 "Straight Waveguide" sch_x=253 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13176 N$26351 N$26352 "Straight Waveguide" sch_x=253 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13177 N$26353 N$26354 "Straight Waveguide" sch_x=253 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13178 N$26355 N$26356 "Straight Waveguide" sch_x=253 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13179 N$26357 N$26358 "Straight Waveguide" sch_x=253 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13180 N$26359 N$26360 "Straight Waveguide" sch_x=253 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13181 N$26361 N$26362 "Straight Waveguide" sch_x=253 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13182 N$26363 N$26364 "Straight Waveguide" sch_x=253 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13183 N$26365 N$26366 "Straight Waveguide" sch_x=253 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13184 N$26367 N$26368 "Straight Waveguide" sch_x=253 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13185 N$26369 N$26370 "Straight Waveguide" sch_x=253 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13186 N$26371 N$26372 "Straight Waveguide" sch_x=253 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13187 N$26373 N$26374 "Straight Waveguide" sch_x=253 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13188 N$26375 N$26376 "Straight Waveguide" sch_x=253 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13189 N$26377 N$26378 "Straight Waveguide" sch_x=253 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13190 N$26379 N$26380 "Straight Waveguide" sch_x=253 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13191 N$26381 N$26382 "Straight Waveguide" sch_x=253 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13192 N$26383 N$26384 "Straight Waveguide" sch_x=253 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13193 N$26385 N$26386 "Straight Waveguide" sch_x=253 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13194 N$26387 N$26388 "Straight Waveguide" sch_x=253 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13195 N$26389 N$26390 "Straight Waveguide" sch_x=253 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13196 N$26391 N$26392 "Straight Waveguide" sch_x=253 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13197 N$26393 N$26394 "Straight Waveguide" sch_x=253 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13198 N$26395 N$26396 "Straight Waveguide" sch_x=253 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13199 N$26397 N$26398 "Straight Waveguide" sch_x=253 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13200 N$26399 N$26400 "Straight Waveguide" sch_x=253 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13201 N$26401 N$26402 "Straight Waveguide" sch_x=253 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13202 N$26403 N$26404 "Straight Waveguide" sch_x=253 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13203 N$26405 N$26406 "Straight Waveguide" sch_x=253 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13204 N$26407 N$26408 "Straight Waveguide" sch_x=253 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13205 N$26409 N$26410 "Straight Waveguide" sch_x=253 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13206 N$26411 N$26412 "Straight Waveguide" sch_x=253 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13207 N$26413 N$26414 "Straight Waveguide" sch_x=253 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13208 N$26415 N$26416 "Straight Waveguide" sch_x=253 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13209 N$26417 N$26418 "Straight Waveguide" sch_x=253 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13210 N$26419 N$26420 "Straight Waveguide" sch_x=253 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13211 N$26421 N$26422 "Straight Waveguide" sch_x=253 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13212 N$26423 N$26424 "Straight Waveguide" sch_x=253 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13213 N$26425 N$26426 "Straight Waveguide" sch_x=253 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13214 N$26427 N$26428 "Straight Waveguide" sch_x=253 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13215 N$26429 N$26430 "Straight Waveguide" sch_x=253 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13216 N$26431 N$26432 "Straight Waveguide" sch_x=253 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13217 N$26433 N$26434 "Straight Waveguide" sch_x=253 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13218 N$26435 N$26436 "Straight Waveguide" sch_x=253 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13219 N$26437 N$26438 "Straight Waveguide" sch_x=253 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13220 N$26439 N$26440 "Straight Waveguide" sch_x=253 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13221 N$26441 N$26442 "Straight Waveguide" sch_x=253 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13222 N$26443 N$26444 "Straight Waveguide" sch_x=253 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13223 N$26445 N$26446 "Straight Waveguide" sch_x=253 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13224 N$26447 N$26448 "Straight Waveguide" sch_x=253 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13225 N$26449 N$26450 "Straight Waveguide" sch_x=253 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13226 N$26451 N$26452 "Straight Waveguide" sch_x=253 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13227 N$26453 N$26454 "Straight Waveguide" sch_x=253 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13228 N$26455 N$26456 "Straight Waveguide" sch_x=253 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13229 N$26457 N$26458 "Straight Waveguide" sch_x=253 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13230 N$26459 N$26460 "Straight Waveguide" sch_x=253 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13231 N$26461 N$26462 "Straight Waveguide" sch_x=253 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13232 N$26463 N$26464 "Straight Waveguide" sch_x=253 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13233 N$26465 N$26466 "Straight Waveguide" sch_x=253 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13234 N$26467 N$26468 "Straight Waveguide" sch_x=253 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13235 N$26469 N$26470 "Straight Waveguide" sch_x=253 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13236 N$26471 N$26472 "Straight Waveguide" sch_x=253 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13237 N$26473 N$26474 "Straight Waveguide" sch_x=253 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13238 N$26475 N$26476 "Straight Waveguide" sch_x=253 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13239 N$26477 N$26478 "Straight Waveguide" sch_x=253 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13240 N$26479 N$26480 "Straight Waveguide" sch_x=253 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13241 N$26481 N$26482 "Straight Waveguide" sch_x=253 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13242 N$26483 N$26484 "Straight Waveguide" sch_x=253 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13243 N$26485 N$26486 "Straight Waveguide" sch_x=253 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13244 N$26487 N$26488 "Straight Waveguide" sch_x=253 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13245 N$26489 N$26490 "Straight Waveguide" sch_x=253 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13246 N$26491 N$26492 "Straight Waveguide" sch_x=253 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13247 N$26493 N$26494 "Straight Waveguide" sch_x=251 sch_y=61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13248 N$26495 N$26496 "Straight Waveguide" sch_x=251 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13249 N$26497 N$26498 "Straight Waveguide" sch_x=251 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13250 N$26499 N$26500 "Straight Waveguide" sch_x=251 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13251 N$26501 N$26502 "Straight Waveguide" sch_x=251 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13252 N$26503 N$26504 "Straight Waveguide" sch_x=251 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13253 N$26505 N$26506 "Straight Waveguide" sch_x=251 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13254 N$26507 N$26508 "Straight Waveguide" sch_x=251 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13255 N$26509 N$26510 "Straight Waveguide" sch_x=251 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13256 N$26511 N$26512 "Straight Waveguide" sch_x=251 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13257 N$26513 N$26514 "Straight Waveguide" sch_x=251 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13258 N$26515 N$26516 "Straight Waveguide" sch_x=251 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13259 N$26517 N$26518 "Straight Waveguide" sch_x=251 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13260 N$26519 N$26520 "Straight Waveguide" sch_x=251 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13261 N$26521 N$26522 "Straight Waveguide" sch_x=251 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13262 N$26523 N$26524 "Straight Waveguide" sch_x=251 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13263 N$26525 N$26526 "Straight Waveguide" sch_x=251 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13264 N$26527 N$26528 "Straight Waveguide" sch_x=251 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13265 N$26529 N$26530 "Straight Waveguide" sch_x=251 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13266 N$26531 N$26532 "Straight Waveguide" sch_x=251 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13267 N$26533 N$26534 "Straight Waveguide" sch_x=251 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13268 N$26535 N$26536 "Straight Waveguide" sch_x=251 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13269 N$26537 N$26538 "Straight Waveguide" sch_x=251 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13270 N$26539 N$26540 "Straight Waveguide" sch_x=251 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13271 N$26541 N$26542 "Straight Waveguide" sch_x=251 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13272 N$26543 N$26544 "Straight Waveguide" sch_x=251 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13273 N$26545 N$26546 "Straight Waveguide" sch_x=251 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13274 N$26547 N$26548 "Straight Waveguide" sch_x=251 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13275 N$26549 N$26550 "Straight Waveguide" sch_x=251 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13276 N$26551 N$26552 "Straight Waveguide" sch_x=251 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13277 N$26553 N$26554 "Straight Waveguide" sch_x=251 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13278 N$26555 N$26556 "Straight Waveguide" sch_x=251 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13279 N$26557 N$26558 "Straight Waveguide" sch_x=251 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13280 N$26559 N$26560 "Straight Waveguide" sch_x=251 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13281 N$26561 N$26562 "Straight Waveguide" sch_x=251 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13282 N$26563 N$26564 "Straight Waveguide" sch_x=251 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13283 N$26565 N$26566 "Straight Waveguide" sch_x=251 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13284 N$26567 N$26568 "Straight Waveguide" sch_x=251 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13285 N$26569 N$26570 "Straight Waveguide" sch_x=251 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13286 N$26571 N$26572 "Straight Waveguide" sch_x=251 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13287 N$26573 N$26574 "Straight Waveguide" sch_x=251 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13288 N$26575 N$26576 "Straight Waveguide" sch_x=251 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13289 N$26577 N$26578 "Straight Waveguide" sch_x=251 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13290 N$26579 N$26580 "Straight Waveguide" sch_x=251 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13291 N$26581 N$26582 "Straight Waveguide" sch_x=251 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13292 N$26583 N$26584 "Straight Waveguide" sch_x=251 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13293 N$26585 N$26586 "Straight Waveguide" sch_x=251 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13294 N$26587 N$26588 "Straight Waveguide" sch_x=251 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13295 N$26589 N$26590 "Straight Waveguide" sch_x=251 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13296 N$26591 N$26592 "Straight Waveguide" sch_x=251 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13297 N$26593 N$26594 "Straight Waveguide" sch_x=251 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13298 N$26595 N$26596 "Straight Waveguide" sch_x=251 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13299 N$26597 N$26598 "Straight Waveguide" sch_x=251 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13300 N$26599 N$26600 "Straight Waveguide" sch_x=251 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13301 N$26601 N$26602 "Straight Waveguide" sch_x=251 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13302 N$26603 N$26604 "Straight Waveguide" sch_x=251 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13303 N$26605 N$26606 "Straight Waveguide" sch_x=251 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13304 N$26607 N$26608 "Straight Waveguide" sch_x=251 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13305 N$26609 N$26610 "Straight Waveguide" sch_x=251 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13306 N$26611 N$26612 "Straight Waveguide" sch_x=251 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13307 N$26613 N$26614 "Straight Waveguide" sch_x=251 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13308 N$26615 N$26616 "Straight Waveguide" sch_x=251 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13309 N$26617 N$26618 "Straight Waveguide" sch_x=251 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13310 N$26619 N$26620 "Straight Waveguide" sch_x=251 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13311 N$26621 N$26622 "Straight Waveguide" sch_x=251 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13312 N$26623 N$26624 "Straight Waveguide" sch_x=251 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13313 N$26625 N$26626 "Straight Waveguide" sch_x=251 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13314 N$26627 N$26628 "Straight Waveguide" sch_x=251 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13315 N$26629 N$26630 "Straight Waveguide" sch_x=251 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13316 N$26631 N$26632 "Straight Waveguide" sch_x=251 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13317 N$26633 N$26634 "Straight Waveguide" sch_x=251 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13318 N$26635 N$26636 "Straight Waveguide" sch_x=251 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13319 N$26637 N$26638 "Straight Waveguide" sch_x=251 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13320 N$26639 N$26640 "Straight Waveguide" sch_x=251 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13321 N$26641 N$26642 "Straight Waveguide" sch_x=251 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13322 N$26643 N$26644 "Straight Waveguide" sch_x=251 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13323 N$26645 N$26646 "Straight Waveguide" sch_x=251 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13324 N$26647 N$26648 "Straight Waveguide" sch_x=251 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13325 N$26649 N$26650 "Straight Waveguide" sch_x=251 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13326 N$26651 N$26652 "Straight Waveguide" sch_x=251 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13327 N$26653 N$26654 "Straight Waveguide" sch_x=251 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13328 N$26655 N$26656 "Straight Waveguide" sch_x=251 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13329 N$26657 N$26658 "Straight Waveguide" sch_x=251 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13330 N$26659 N$26660 "Straight Waveguide" sch_x=251 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13331 N$26661 N$26662 "Straight Waveguide" sch_x=251 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13332 N$26663 N$26664 "Straight Waveguide" sch_x=251 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13333 N$26665 N$26666 "Straight Waveguide" sch_x=251 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13334 N$26667 N$26668 "Straight Waveguide" sch_x=251 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13335 N$26669 N$26670 "Straight Waveguide" sch_x=251 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13336 N$26671 N$26672 "Straight Waveguide" sch_x=251 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13337 N$26673 N$26674 "Straight Waveguide" sch_x=251 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13338 N$26675 N$26676 "Straight Waveguide" sch_x=251 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13339 N$26677 N$26678 "Straight Waveguide" sch_x=251 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13340 N$26679 N$26680 "Straight Waveguide" sch_x=251 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13341 N$26681 N$26682 "Straight Waveguide" sch_x=251 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13342 N$26683 N$26684 "Straight Waveguide" sch_x=251 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13343 N$26685 N$26686 "Straight Waveguide" sch_x=251 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13344 N$26687 N$26688 "Straight Waveguide" sch_x=251 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13345 N$26689 N$26690 "Straight Waveguide" sch_x=251 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13346 N$26691 N$26692 "Straight Waveguide" sch_x=251 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13347 N$26693 N$26694 "Straight Waveguide" sch_x=251 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13348 N$26695 N$26696 "Straight Waveguide" sch_x=251 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13349 N$26697 N$26698 "Straight Waveguide" sch_x=251 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13350 N$26699 N$26700 "Straight Waveguide" sch_x=251 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13351 N$26701 N$26702 "Straight Waveguide" sch_x=251 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13352 N$26703 N$26704 "Straight Waveguide" sch_x=251 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13353 N$26705 N$26706 "Straight Waveguide" sch_x=251 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13354 N$26707 N$26708 "Straight Waveguide" sch_x=251 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13355 N$26709 N$26710 "Straight Waveguide" sch_x=251 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13356 N$26711 N$26712 "Straight Waveguide" sch_x=251 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13357 N$26713 N$26714 "Straight Waveguide" sch_x=251 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13358 N$26715 N$26716 "Straight Waveguide" sch_x=251 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13359 N$26717 N$26718 "Straight Waveguide" sch_x=251 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13360 N$26719 N$26720 "Straight Waveguide" sch_x=251 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13361 N$26721 N$26722 "Straight Waveguide" sch_x=251 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13362 N$26723 N$26724 "Straight Waveguide" sch_x=251 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13363 N$26725 N$26726 "Straight Waveguide" sch_x=251 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13364 N$26727 N$26728 "Straight Waveguide" sch_x=251 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13365 N$26729 N$26730 "Straight Waveguide" sch_x=251 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13366 N$26731 N$26732 "Straight Waveguide" sch_x=251 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13367 N$26733 N$26734 "Straight Waveguide" sch_x=251 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13368 N$26735 N$26736 "Straight Waveguide" sch_x=251 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13369 N$26737 N$26738 "Straight Waveguide" sch_x=251 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13370 N$26739 N$26740 "Straight Waveguide" sch_x=251 sch_y=-61.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13371 N$26741 N$26742 "Straight Waveguide" sch_x=249 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13372 N$26743 N$26744 "Straight Waveguide" sch_x=249 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13373 N$26745 N$26746 "Straight Waveguide" sch_x=249 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13374 N$26747 N$26748 "Straight Waveguide" sch_x=249 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13375 N$26749 N$26750 "Straight Waveguide" sch_x=249 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13376 N$26751 N$26752 "Straight Waveguide" sch_x=249 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13377 N$26753 N$26754 "Straight Waveguide" sch_x=249 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13378 N$26755 N$26756 "Straight Waveguide" sch_x=249 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13379 N$26757 N$26758 "Straight Waveguide" sch_x=249 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13380 N$26759 N$26760 "Straight Waveguide" sch_x=249 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13381 N$26761 N$26762 "Straight Waveguide" sch_x=249 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13382 N$26763 N$26764 "Straight Waveguide" sch_x=249 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13383 N$26765 N$26766 "Straight Waveguide" sch_x=249 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13384 N$26767 N$26768 "Straight Waveguide" sch_x=249 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13385 N$26769 N$26770 "Straight Waveguide" sch_x=249 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13386 N$26771 N$26772 "Straight Waveguide" sch_x=249 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13387 N$26773 N$26774 "Straight Waveguide" sch_x=249 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13388 N$26775 N$26776 "Straight Waveguide" sch_x=249 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13389 N$26777 N$26778 "Straight Waveguide" sch_x=249 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13390 N$26779 N$26780 "Straight Waveguide" sch_x=249 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13391 N$26781 N$26782 "Straight Waveguide" sch_x=249 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13392 N$26783 N$26784 "Straight Waveguide" sch_x=249 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13393 N$26785 N$26786 "Straight Waveguide" sch_x=249 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13394 N$26787 N$26788 "Straight Waveguide" sch_x=249 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13395 N$26789 N$26790 "Straight Waveguide" sch_x=249 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13396 N$26791 N$26792 "Straight Waveguide" sch_x=249 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13397 N$26793 N$26794 "Straight Waveguide" sch_x=249 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13398 N$26795 N$26796 "Straight Waveguide" sch_x=249 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13399 N$26797 N$26798 "Straight Waveguide" sch_x=249 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13400 N$26799 N$26800 "Straight Waveguide" sch_x=249 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13401 N$26801 N$26802 "Straight Waveguide" sch_x=249 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13402 N$26803 N$26804 "Straight Waveguide" sch_x=249 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13403 N$26805 N$26806 "Straight Waveguide" sch_x=249 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13404 N$26807 N$26808 "Straight Waveguide" sch_x=249 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13405 N$26809 N$26810 "Straight Waveguide" sch_x=249 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13406 N$26811 N$26812 "Straight Waveguide" sch_x=249 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13407 N$26813 N$26814 "Straight Waveguide" sch_x=249 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13408 N$26815 N$26816 "Straight Waveguide" sch_x=249 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13409 N$26817 N$26818 "Straight Waveguide" sch_x=249 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13410 N$26819 N$26820 "Straight Waveguide" sch_x=249 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13411 N$26821 N$26822 "Straight Waveguide" sch_x=249 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13412 N$26823 N$26824 "Straight Waveguide" sch_x=249 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13413 N$26825 N$26826 "Straight Waveguide" sch_x=249 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13414 N$26827 N$26828 "Straight Waveguide" sch_x=249 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13415 N$26829 N$26830 "Straight Waveguide" sch_x=249 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13416 N$26831 N$26832 "Straight Waveguide" sch_x=249 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13417 N$26833 N$26834 "Straight Waveguide" sch_x=249 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13418 N$26835 N$26836 "Straight Waveguide" sch_x=249 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13419 N$26837 N$26838 "Straight Waveguide" sch_x=249 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13420 N$26839 N$26840 "Straight Waveguide" sch_x=249 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13421 N$26841 N$26842 "Straight Waveguide" sch_x=249 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13422 N$26843 N$26844 "Straight Waveguide" sch_x=249 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13423 N$26845 N$26846 "Straight Waveguide" sch_x=249 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13424 N$26847 N$26848 "Straight Waveguide" sch_x=249 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13425 N$26849 N$26850 "Straight Waveguide" sch_x=249 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13426 N$26851 N$26852 "Straight Waveguide" sch_x=249 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13427 N$26853 N$26854 "Straight Waveguide" sch_x=249 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13428 N$26855 N$26856 "Straight Waveguide" sch_x=249 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13429 N$26857 N$26858 "Straight Waveguide" sch_x=249 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13430 N$26859 N$26860 "Straight Waveguide" sch_x=249 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13431 N$26861 N$26862 "Straight Waveguide" sch_x=249 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13432 N$26863 N$26864 "Straight Waveguide" sch_x=249 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13433 N$26865 N$26866 "Straight Waveguide" sch_x=249 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13434 N$26867 N$26868 "Straight Waveguide" sch_x=249 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13435 N$26869 N$26870 "Straight Waveguide" sch_x=249 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13436 N$26871 N$26872 "Straight Waveguide" sch_x=249 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13437 N$26873 N$26874 "Straight Waveguide" sch_x=249 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13438 N$26875 N$26876 "Straight Waveguide" sch_x=249 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13439 N$26877 N$26878 "Straight Waveguide" sch_x=249 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13440 N$26879 N$26880 "Straight Waveguide" sch_x=249 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13441 N$26881 N$26882 "Straight Waveguide" sch_x=249 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13442 N$26883 N$26884 "Straight Waveguide" sch_x=249 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13443 N$26885 N$26886 "Straight Waveguide" sch_x=249 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13444 N$26887 N$26888 "Straight Waveguide" sch_x=249 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13445 N$26889 N$26890 "Straight Waveguide" sch_x=249 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13446 N$26891 N$26892 "Straight Waveguide" sch_x=249 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13447 N$26893 N$26894 "Straight Waveguide" sch_x=249 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13448 N$26895 N$26896 "Straight Waveguide" sch_x=249 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13449 N$26897 N$26898 "Straight Waveguide" sch_x=249 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13450 N$26899 N$26900 "Straight Waveguide" sch_x=249 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13451 N$26901 N$26902 "Straight Waveguide" sch_x=249 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13452 N$26903 N$26904 "Straight Waveguide" sch_x=249 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13453 N$26905 N$26906 "Straight Waveguide" sch_x=249 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13454 N$26907 N$26908 "Straight Waveguide" sch_x=249 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13455 N$26909 N$26910 "Straight Waveguide" sch_x=249 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13456 N$26911 N$26912 "Straight Waveguide" sch_x=249 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13457 N$26913 N$26914 "Straight Waveguide" sch_x=249 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13458 N$26915 N$26916 "Straight Waveguide" sch_x=249 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13459 N$26917 N$26918 "Straight Waveguide" sch_x=249 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13460 N$26919 N$26920 "Straight Waveguide" sch_x=249 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13461 N$26921 N$26922 "Straight Waveguide" sch_x=249 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13462 N$26923 N$26924 "Straight Waveguide" sch_x=249 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13463 N$26925 N$26926 "Straight Waveguide" sch_x=249 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13464 N$26927 N$26928 "Straight Waveguide" sch_x=249 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13465 N$26929 N$26930 "Straight Waveguide" sch_x=249 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13466 N$26931 N$26932 "Straight Waveguide" sch_x=249 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13467 N$26933 N$26934 "Straight Waveguide" sch_x=249 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13468 N$26935 N$26936 "Straight Waveguide" sch_x=249 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13469 N$26937 N$26938 "Straight Waveguide" sch_x=249 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13470 N$26939 N$26940 "Straight Waveguide" sch_x=249 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13471 N$26941 N$26942 "Straight Waveguide" sch_x=249 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13472 N$26943 N$26944 "Straight Waveguide" sch_x=249 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13473 N$26945 N$26946 "Straight Waveguide" sch_x=249 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13474 N$26947 N$26948 "Straight Waveguide" sch_x=249 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13475 N$26949 N$26950 "Straight Waveguide" sch_x=249 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13476 N$26951 N$26952 "Straight Waveguide" sch_x=249 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13477 N$26953 N$26954 "Straight Waveguide" sch_x=249 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13478 N$26955 N$26956 "Straight Waveguide" sch_x=249 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13479 N$26957 N$26958 "Straight Waveguide" sch_x=249 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13480 N$26959 N$26960 "Straight Waveguide" sch_x=249 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13481 N$26961 N$26962 "Straight Waveguide" sch_x=249 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13482 N$26963 N$26964 "Straight Waveguide" sch_x=249 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13483 N$26965 N$26966 "Straight Waveguide" sch_x=249 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13484 N$26967 N$26968 "Straight Waveguide" sch_x=249 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13485 N$26969 N$26970 "Straight Waveguide" sch_x=249 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13486 N$26971 N$26972 "Straight Waveguide" sch_x=249 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13487 N$26973 N$26974 "Straight Waveguide" sch_x=249 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13488 N$26975 N$26976 "Straight Waveguide" sch_x=249 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13489 N$26977 N$26978 "Straight Waveguide" sch_x=249 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13490 N$26979 N$26980 "Straight Waveguide" sch_x=249 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13491 N$26981 N$26982 "Straight Waveguide" sch_x=249 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13492 N$26983 N$26984 "Straight Waveguide" sch_x=249 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13493 N$26985 N$26986 "Straight Waveguide" sch_x=247 sch_y=59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13494 N$26987 N$26988 "Straight Waveguide" sch_x=247 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13495 N$26989 N$26990 "Straight Waveguide" sch_x=247 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13496 N$26991 N$26992 "Straight Waveguide" sch_x=247 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13497 N$26993 N$26994 "Straight Waveguide" sch_x=247 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13498 N$26995 N$26996 "Straight Waveguide" sch_x=247 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13499 N$26997 N$26998 "Straight Waveguide" sch_x=247 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13500 N$26999 N$27000 "Straight Waveguide" sch_x=247 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13501 N$27001 N$27002 "Straight Waveguide" sch_x=247 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13502 N$27003 N$27004 "Straight Waveguide" sch_x=247 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13503 N$27005 N$27006 "Straight Waveguide" sch_x=247 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13504 N$27007 N$27008 "Straight Waveguide" sch_x=247 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13505 N$27009 N$27010 "Straight Waveguide" sch_x=247 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13506 N$27011 N$27012 "Straight Waveguide" sch_x=247 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13507 N$27013 N$27014 "Straight Waveguide" sch_x=247 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13508 N$27015 N$27016 "Straight Waveguide" sch_x=247 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13509 N$27017 N$27018 "Straight Waveguide" sch_x=247 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13510 N$27019 N$27020 "Straight Waveguide" sch_x=247 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13511 N$27021 N$27022 "Straight Waveguide" sch_x=247 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13512 N$27023 N$27024 "Straight Waveguide" sch_x=247 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13513 N$27025 N$27026 "Straight Waveguide" sch_x=247 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13514 N$27027 N$27028 "Straight Waveguide" sch_x=247 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13515 N$27029 N$27030 "Straight Waveguide" sch_x=247 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13516 N$27031 N$27032 "Straight Waveguide" sch_x=247 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13517 N$27033 N$27034 "Straight Waveguide" sch_x=247 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13518 N$27035 N$27036 "Straight Waveguide" sch_x=247 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13519 N$27037 N$27038 "Straight Waveguide" sch_x=247 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13520 N$27039 N$27040 "Straight Waveguide" sch_x=247 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13521 N$27041 N$27042 "Straight Waveguide" sch_x=247 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13522 N$27043 N$27044 "Straight Waveguide" sch_x=247 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13523 N$27045 N$27046 "Straight Waveguide" sch_x=247 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13524 N$27047 N$27048 "Straight Waveguide" sch_x=247 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13525 N$27049 N$27050 "Straight Waveguide" sch_x=247 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13526 N$27051 N$27052 "Straight Waveguide" sch_x=247 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13527 N$27053 N$27054 "Straight Waveguide" sch_x=247 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13528 N$27055 N$27056 "Straight Waveguide" sch_x=247 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13529 N$27057 N$27058 "Straight Waveguide" sch_x=247 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13530 N$27059 N$27060 "Straight Waveguide" sch_x=247 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13531 N$27061 N$27062 "Straight Waveguide" sch_x=247 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13532 N$27063 N$27064 "Straight Waveguide" sch_x=247 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13533 N$27065 N$27066 "Straight Waveguide" sch_x=247 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13534 N$27067 N$27068 "Straight Waveguide" sch_x=247 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13535 N$27069 N$27070 "Straight Waveguide" sch_x=247 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13536 N$27071 N$27072 "Straight Waveguide" sch_x=247 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13537 N$27073 N$27074 "Straight Waveguide" sch_x=247 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13538 N$27075 N$27076 "Straight Waveguide" sch_x=247 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13539 N$27077 N$27078 "Straight Waveguide" sch_x=247 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13540 N$27079 N$27080 "Straight Waveguide" sch_x=247 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13541 N$27081 N$27082 "Straight Waveguide" sch_x=247 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13542 N$27083 N$27084 "Straight Waveguide" sch_x=247 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13543 N$27085 N$27086 "Straight Waveguide" sch_x=247 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13544 N$27087 N$27088 "Straight Waveguide" sch_x=247 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13545 N$27089 N$27090 "Straight Waveguide" sch_x=247 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13546 N$27091 N$27092 "Straight Waveguide" sch_x=247 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13547 N$27093 N$27094 "Straight Waveguide" sch_x=247 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13548 N$27095 N$27096 "Straight Waveguide" sch_x=247 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13549 N$27097 N$27098 "Straight Waveguide" sch_x=247 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13550 N$27099 N$27100 "Straight Waveguide" sch_x=247 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13551 N$27101 N$27102 "Straight Waveguide" sch_x=247 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13552 N$27103 N$27104 "Straight Waveguide" sch_x=247 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13553 N$27105 N$27106 "Straight Waveguide" sch_x=247 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13554 N$27107 N$27108 "Straight Waveguide" sch_x=247 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13555 N$27109 N$27110 "Straight Waveguide" sch_x=247 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13556 N$27111 N$27112 "Straight Waveguide" sch_x=247 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13557 N$27113 N$27114 "Straight Waveguide" sch_x=247 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13558 N$27115 N$27116 "Straight Waveguide" sch_x=247 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13559 N$27117 N$27118 "Straight Waveguide" sch_x=247 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13560 N$27119 N$27120 "Straight Waveguide" sch_x=247 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13561 N$27121 N$27122 "Straight Waveguide" sch_x=247 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13562 N$27123 N$27124 "Straight Waveguide" sch_x=247 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13563 N$27125 N$27126 "Straight Waveguide" sch_x=247 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13564 N$27127 N$27128 "Straight Waveguide" sch_x=247 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13565 N$27129 N$27130 "Straight Waveguide" sch_x=247 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13566 N$27131 N$27132 "Straight Waveguide" sch_x=247 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13567 N$27133 N$27134 "Straight Waveguide" sch_x=247 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13568 N$27135 N$27136 "Straight Waveguide" sch_x=247 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13569 N$27137 N$27138 "Straight Waveguide" sch_x=247 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13570 N$27139 N$27140 "Straight Waveguide" sch_x=247 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13571 N$27141 N$27142 "Straight Waveguide" sch_x=247 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13572 N$27143 N$27144 "Straight Waveguide" sch_x=247 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13573 N$27145 N$27146 "Straight Waveguide" sch_x=247 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13574 N$27147 N$27148 "Straight Waveguide" sch_x=247 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13575 N$27149 N$27150 "Straight Waveguide" sch_x=247 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13576 N$27151 N$27152 "Straight Waveguide" sch_x=247 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13577 N$27153 N$27154 "Straight Waveguide" sch_x=247 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13578 N$27155 N$27156 "Straight Waveguide" sch_x=247 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13579 N$27157 N$27158 "Straight Waveguide" sch_x=247 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13580 N$27159 N$27160 "Straight Waveguide" sch_x=247 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13581 N$27161 N$27162 "Straight Waveguide" sch_x=247 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13582 N$27163 N$27164 "Straight Waveguide" sch_x=247 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13583 N$27165 N$27166 "Straight Waveguide" sch_x=247 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13584 N$27167 N$27168 "Straight Waveguide" sch_x=247 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13585 N$27169 N$27170 "Straight Waveguide" sch_x=247 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13586 N$27171 N$27172 "Straight Waveguide" sch_x=247 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13587 N$27173 N$27174 "Straight Waveguide" sch_x=247 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13588 N$27175 N$27176 "Straight Waveguide" sch_x=247 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13589 N$27177 N$27178 "Straight Waveguide" sch_x=247 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13590 N$27179 N$27180 "Straight Waveguide" sch_x=247 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13591 N$27181 N$27182 "Straight Waveguide" sch_x=247 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13592 N$27183 N$27184 "Straight Waveguide" sch_x=247 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13593 N$27185 N$27186 "Straight Waveguide" sch_x=247 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13594 N$27187 N$27188 "Straight Waveguide" sch_x=247 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13595 N$27189 N$27190 "Straight Waveguide" sch_x=247 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13596 N$27191 N$27192 "Straight Waveguide" sch_x=247 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13597 N$27193 N$27194 "Straight Waveguide" sch_x=247 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13598 N$27195 N$27196 "Straight Waveguide" sch_x=247 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13599 N$27197 N$27198 "Straight Waveguide" sch_x=247 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13600 N$27199 N$27200 "Straight Waveguide" sch_x=247 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13601 N$27201 N$27202 "Straight Waveguide" sch_x=247 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13602 N$27203 N$27204 "Straight Waveguide" sch_x=247 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13603 N$27205 N$27206 "Straight Waveguide" sch_x=247 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13604 N$27207 N$27208 "Straight Waveguide" sch_x=247 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13605 N$27209 N$27210 "Straight Waveguide" sch_x=247 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13606 N$27211 N$27212 "Straight Waveguide" sch_x=247 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13607 N$27213 N$27214 "Straight Waveguide" sch_x=247 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13608 N$27215 N$27216 "Straight Waveguide" sch_x=247 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13609 N$27217 N$27218 "Straight Waveguide" sch_x=247 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13610 N$27219 N$27220 "Straight Waveguide" sch_x=247 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13611 N$27221 N$27222 "Straight Waveguide" sch_x=247 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13612 N$27223 N$27224 "Straight Waveguide" sch_x=247 sch_y=-59.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13613 N$27225 N$27226 "Straight Waveguide" sch_x=245 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13614 N$27227 N$27228 "Straight Waveguide" sch_x=245 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13615 N$27229 N$27230 "Straight Waveguide" sch_x=245 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13616 N$27231 N$27232 "Straight Waveguide" sch_x=245 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13617 N$27233 N$27234 "Straight Waveguide" sch_x=245 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13618 N$27235 N$27236 "Straight Waveguide" sch_x=245 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13619 N$27237 N$27238 "Straight Waveguide" sch_x=245 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13620 N$27239 N$27240 "Straight Waveguide" sch_x=245 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13621 N$27241 N$27242 "Straight Waveguide" sch_x=245 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13622 N$27243 N$27244 "Straight Waveguide" sch_x=245 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13623 N$27245 N$27246 "Straight Waveguide" sch_x=245 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13624 N$27247 N$27248 "Straight Waveguide" sch_x=245 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13625 N$27249 N$27250 "Straight Waveguide" sch_x=245 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13626 N$27251 N$27252 "Straight Waveguide" sch_x=245 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13627 N$27253 N$27254 "Straight Waveguide" sch_x=245 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13628 N$27255 N$27256 "Straight Waveguide" sch_x=245 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13629 N$27257 N$27258 "Straight Waveguide" sch_x=245 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13630 N$27259 N$27260 "Straight Waveguide" sch_x=245 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13631 N$27261 N$27262 "Straight Waveguide" sch_x=245 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13632 N$27263 N$27264 "Straight Waveguide" sch_x=245 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13633 N$27265 N$27266 "Straight Waveguide" sch_x=245 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13634 N$27267 N$27268 "Straight Waveguide" sch_x=245 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13635 N$27269 N$27270 "Straight Waveguide" sch_x=245 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13636 N$27271 N$27272 "Straight Waveguide" sch_x=245 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13637 N$27273 N$27274 "Straight Waveguide" sch_x=245 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13638 N$27275 N$27276 "Straight Waveguide" sch_x=245 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13639 N$27277 N$27278 "Straight Waveguide" sch_x=245 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13640 N$27279 N$27280 "Straight Waveguide" sch_x=245 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13641 N$27281 N$27282 "Straight Waveguide" sch_x=245 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13642 N$27283 N$27284 "Straight Waveguide" sch_x=245 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13643 N$27285 N$27286 "Straight Waveguide" sch_x=245 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13644 N$27287 N$27288 "Straight Waveguide" sch_x=245 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13645 N$27289 N$27290 "Straight Waveguide" sch_x=245 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13646 N$27291 N$27292 "Straight Waveguide" sch_x=245 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13647 N$27293 N$27294 "Straight Waveguide" sch_x=245 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13648 N$27295 N$27296 "Straight Waveguide" sch_x=245 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13649 N$27297 N$27298 "Straight Waveguide" sch_x=245 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13650 N$27299 N$27300 "Straight Waveguide" sch_x=245 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13651 N$27301 N$27302 "Straight Waveguide" sch_x=245 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13652 N$27303 N$27304 "Straight Waveguide" sch_x=245 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13653 N$27305 N$27306 "Straight Waveguide" sch_x=245 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13654 N$27307 N$27308 "Straight Waveguide" sch_x=245 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13655 N$27309 N$27310 "Straight Waveguide" sch_x=245 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13656 N$27311 N$27312 "Straight Waveguide" sch_x=245 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13657 N$27313 N$27314 "Straight Waveguide" sch_x=245 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13658 N$27315 N$27316 "Straight Waveguide" sch_x=245 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13659 N$27317 N$27318 "Straight Waveguide" sch_x=245 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13660 N$27319 N$27320 "Straight Waveguide" sch_x=245 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13661 N$27321 N$27322 "Straight Waveguide" sch_x=245 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13662 N$27323 N$27324 "Straight Waveguide" sch_x=245 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13663 N$27325 N$27326 "Straight Waveguide" sch_x=245 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13664 N$27327 N$27328 "Straight Waveguide" sch_x=245 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13665 N$27329 N$27330 "Straight Waveguide" sch_x=245 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13666 N$27331 N$27332 "Straight Waveguide" sch_x=245 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13667 N$27333 N$27334 "Straight Waveguide" sch_x=245 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13668 N$27335 N$27336 "Straight Waveguide" sch_x=245 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13669 N$27337 N$27338 "Straight Waveguide" sch_x=245 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13670 N$27339 N$27340 "Straight Waveguide" sch_x=245 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13671 N$27341 N$27342 "Straight Waveguide" sch_x=245 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13672 N$27343 N$27344 "Straight Waveguide" sch_x=245 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13673 N$27345 N$27346 "Straight Waveguide" sch_x=245 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13674 N$27347 N$27348 "Straight Waveguide" sch_x=245 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13675 N$27349 N$27350 "Straight Waveguide" sch_x=245 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13676 N$27351 N$27352 "Straight Waveguide" sch_x=245 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13677 N$27353 N$27354 "Straight Waveguide" sch_x=245 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13678 N$27355 N$27356 "Straight Waveguide" sch_x=245 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13679 N$27357 N$27358 "Straight Waveguide" sch_x=245 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13680 N$27359 N$27360 "Straight Waveguide" sch_x=245 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13681 N$27361 N$27362 "Straight Waveguide" sch_x=245 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13682 N$27363 N$27364 "Straight Waveguide" sch_x=245 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13683 N$27365 N$27366 "Straight Waveguide" sch_x=245 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13684 N$27367 N$27368 "Straight Waveguide" sch_x=245 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13685 N$27369 N$27370 "Straight Waveguide" sch_x=245 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13686 N$27371 N$27372 "Straight Waveguide" sch_x=245 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13687 N$27373 N$27374 "Straight Waveguide" sch_x=245 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13688 N$27375 N$27376 "Straight Waveguide" sch_x=245 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13689 N$27377 N$27378 "Straight Waveguide" sch_x=245 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13690 N$27379 N$27380 "Straight Waveguide" sch_x=245 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13691 N$27381 N$27382 "Straight Waveguide" sch_x=245 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13692 N$27383 N$27384 "Straight Waveguide" sch_x=245 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13693 N$27385 N$27386 "Straight Waveguide" sch_x=245 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13694 N$27387 N$27388 "Straight Waveguide" sch_x=245 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13695 N$27389 N$27390 "Straight Waveguide" sch_x=245 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13696 N$27391 N$27392 "Straight Waveguide" sch_x=245 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13697 N$27393 N$27394 "Straight Waveguide" sch_x=245 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13698 N$27395 N$27396 "Straight Waveguide" sch_x=245 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13699 N$27397 N$27398 "Straight Waveguide" sch_x=245 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13700 N$27399 N$27400 "Straight Waveguide" sch_x=245 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13701 N$27401 N$27402 "Straight Waveguide" sch_x=245 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13702 N$27403 N$27404 "Straight Waveguide" sch_x=245 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13703 N$27405 N$27406 "Straight Waveguide" sch_x=245 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13704 N$27407 N$27408 "Straight Waveguide" sch_x=245 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13705 N$27409 N$27410 "Straight Waveguide" sch_x=245 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13706 N$27411 N$27412 "Straight Waveguide" sch_x=245 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13707 N$27413 N$27414 "Straight Waveguide" sch_x=245 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13708 N$27415 N$27416 "Straight Waveguide" sch_x=245 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13709 N$27417 N$27418 "Straight Waveguide" sch_x=245 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13710 N$27419 N$27420 "Straight Waveguide" sch_x=245 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13711 N$27421 N$27422 "Straight Waveguide" sch_x=245 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13712 N$27423 N$27424 "Straight Waveguide" sch_x=245 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13713 N$27425 N$27426 "Straight Waveguide" sch_x=245 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13714 N$27427 N$27428 "Straight Waveguide" sch_x=245 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13715 N$27429 N$27430 "Straight Waveguide" sch_x=245 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13716 N$27431 N$27432 "Straight Waveguide" sch_x=245 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13717 N$27433 N$27434 "Straight Waveguide" sch_x=245 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13718 N$27435 N$27436 "Straight Waveguide" sch_x=245 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13719 N$27437 N$27438 "Straight Waveguide" sch_x=245 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13720 N$27439 N$27440 "Straight Waveguide" sch_x=245 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13721 N$27441 N$27442 "Straight Waveguide" sch_x=245 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13722 N$27443 N$27444 "Straight Waveguide" sch_x=245 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13723 N$27445 N$27446 "Straight Waveguide" sch_x=245 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13724 N$27447 N$27448 "Straight Waveguide" sch_x=245 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13725 N$27449 N$27450 "Straight Waveguide" sch_x=245 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13726 N$27451 N$27452 "Straight Waveguide" sch_x=245 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13727 N$27453 N$27454 "Straight Waveguide" sch_x=245 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13728 N$27455 N$27456 "Straight Waveguide" sch_x=245 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13729 N$27457 N$27458 "Straight Waveguide" sch_x=245 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13730 N$27459 N$27460 "Straight Waveguide" sch_x=245 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13731 N$27461 N$27462 "Straight Waveguide" sch_x=243 sch_y=57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13732 N$27463 N$27464 "Straight Waveguide" sch_x=243 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13733 N$27465 N$27466 "Straight Waveguide" sch_x=243 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13734 N$27467 N$27468 "Straight Waveguide" sch_x=243 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13735 N$27469 N$27470 "Straight Waveguide" sch_x=243 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13736 N$27471 N$27472 "Straight Waveguide" sch_x=243 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13737 N$27473 N$27474 "Straight Waveguide" sch_x=243 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13738 N$27475 N$27476 "Straight Waveguide" sch_x=243 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13739 N$27477 N$27478 "Straight Waveguide" sch_x=243 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13740 N$27479 N$27480 "Straight Waveguide" sch_x=243 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13741 N$27481 N$27482 "Straight Waveguide" sch_x=243 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13742 N$27483 N$27484 "Straight Waveguide" sch_x=243 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13743 N$27485 N$27486 "Straight Waveguide" sch_x=243 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13744 N$27487 N$27488 "Straight Waveguide" sch_x=243 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13745 N$27489 N$27490 "Straight Waveguide" sch_x=243 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13746 N$27491 N$27492 "Straight Waveguide" sch_x=243 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13747 N$27493 N$27494 "Straight Waveguide" sch_x=243 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13748 N$27495 N$27496 "Straight Waveguide" sch_x=243 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13749 N$27497 N$27498 "Straight Waveguide" sch_x=243 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13750 N$27499 N$27500 "Straight Waveguide" sch_x=243 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13751 N$27501 N$27502 "Straight Waveguide" sch_x=243 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13752 N$27503 N$27504 "Straight Waveguide" sch_x=243 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13753 N$27505 N$27506 "Straight Waveguide" sch_x=243 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13754 N$27507 N$27508 "Straight Waveguide" sch_x=243 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13755 N$27509 N$27510 "Straight Waveguide" sch_x=243 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13756 N$27511 N$27512 "Straight Waveguide" sch_x=243 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13757 N$27513 N$27514 "Straight Waveguide" sch_x=243 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13758 N$27515 N$27516 "Straight Waveguide" sch_x=243 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13759 N$27517 N$27518 "Straight Waveguide" sch_x=243 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13760 N$27519 N$27520 "Straight Waveguide" sch_x=243 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13761 N$27521 N$27522 "Straight Waveguide" sch_x=243 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13762 N$27523 N$27524 "Straight Waveguide" sch_x=243 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13763 N$27525 N$27526 "Straight Waveguide" sch_x=243 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13764 N$27527 N$27528 "Straight Waveguide" sch_x=243 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13765 N$27529 N$27530 "Straight Waveguide" sch_x=243 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13766 N$27531 N$27532 "Straight Waveguide" sch_x=243 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13767 N$27533 N$27534 "Straight Waveguide" sch_x=243 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13768 N$27535 N$27536 "Straight Waveguide" sch_x=243 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13769 N$27537 N$27538 "Straight Waveguide" sch_x=243 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13770 N$27539 N$27540 "Straight Waveguide" sch_x=243 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13771 N$27541 N$27542 "Straight Waveguide" sch_x=243 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13772 N$27543 N$27544 "Straight Waveguide" sch_x=243 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13773 N$27545 N$27546 "Straight Waveguide" sch_x=243 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13774 N$27547 N$27548 "Straight Waveguide" sch_x=243 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13775 N$27549 N$27550 "Straight Waveguide" sch_x=243 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13776 N$27551 N$27552 "Straight Waveguide" sch_x=243 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13777 N$27553 N$27554 "Straight Waveguide" sch_x=243 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13778 N$27555 N$27556 "Straight Waveguide" sch_x=243 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13779 N$27557 N$27558 "Straight Waveguide" sch_x=243 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13780 N$27559 N$27560 "Straight Waveguide" sch_x=243 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13781 N$27561 N$27562 "Straight Waveguide" sch_x=243 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13782 N$27563 N$27564 "Straight Waveguide" sch_x=243 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13783 N$27565 N$27566 "Straight Waveguide" sch_x=243 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13784 N$27567 N$27568 "Straight Waveguide" sch_x=243 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13785 N$27569 N$27570 "Straight Waveguide" sch_x=243 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13786 N$27571 N$27572 "Straight Waveguide" sch_x=243 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13787 N$27573 N$27574 "Straight Waveguide" sch_x=243 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13788 N$27575 N$27576 "Straight Waveguide" sch_x=243 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13789 N$27577 N$27578 "Straight Waveguide" sch_x=243 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13790 N$27579 N$27580 "Straight Waveguide" sch_x=243 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13791 N$27581 N$27582 "Straight Waveguide" sch_x=243 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13792 N$27583 N$27584 "Straight Waveguide" sch_x=243 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13793 N$27585 N$27586 "Straight Waveguide" sch_x=243 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13794 N$27587 N$27588 "Straight Waveguide" sch_x=243 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13795 N$27589 N$27590 "Straight Waveguide" sch_x=243 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13796 N$27591 N$27592 "Straight Waveguide" sch_x=243 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13797 N$27593 N$27594 "Straight Waveguide" sch_x=243 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13798 N$27595 N$27596 "Straight Waveguide" sch_x=243 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13799 N$27597 N$27598 "Straight Waveguide" sch_x=243 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13800 N$27599 N$27600 "Straight Waveguide" sch_x=243 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13801 N$27601 N$27602 "Straight Waveguide" sch_x=243 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13802 N$27603 N$27604 "Straight Waveguide" sch_x=243 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13803 N$27605 N$27606 "Straight Waveguide" sch_x=243 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13804 N$27607 N$27608 "Straight Waveguide" sch_x=243 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13805 N$27609 N$27610 "Straight Waveguide" sch_x=243 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13806 N$27611 N$27612 "Straight Waveguide" sch_x=243 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13807 N$27613 N$27614 "Straight Waveguide" sch_x=243 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13808 N$27615 N$27616 "Straight Waveguide" sch_x=243 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13809 N$27617 N$27618 "Straight Waveguide" sch_x=243 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13810 N$27619 N$27620 "Straight Waveguide" sch_x=243 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13811 N$27621 N$27622 "Straight Waveguide" sch_x=243 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13812 N$27623 N$27624 "Straight Waveguide" sch_x=243 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13813 N$27625 N$27626 "Straight Waveguide" sch_x=243 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13814 N$27627 N$27628 "Straight Waveguide" sch_x=243 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13815 N$27629 N$27630 "Straight Waveguide" sch_x=243 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13816 N$27631 N$27632 "Straight Waveguide" sch_x=243 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13817 N$27633 N$27634 "Straight Waveguide" sch_x=243 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13818 N$27635 N$27636 "Straight Waveguide" sch_x=243 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13819 N$27637 N$27638 "Straight Waveguide" sch_x=243 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13820 N$27639 N$27640 "Straight Waveguide" sch_x=243 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13821 N$27641 N$27642 "Straight Waveguide" sch_x=243 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13822 N$27643 N$27644 "Straight Waveguide" sch_x=243 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13823 N$27645 N$27646 "Straight Waveguide" sch_x=243 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13824 N$27647 N$27648 "Straight Waveguide" sch_x=243 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13825 N$27649 N$27650 "Straight Waveguide" sch_x=243 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13826 N$27651 N$27652 "Straight Waveguide" sch_x=243 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13827 N$27653 N$27654 "Straight Waveguide" sch_x=243 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13828 N$27655 N$27656 "Straight Waveguide" sch_x=243 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13829 N$27657 N$27658 "Straight Waveguide" sch_x=243 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13830 N$27659 N$27660 "Straight Waveguide" sch_x=243 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13831 N$27661 N$27662 "Straight Waveguide" sch_x=243 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13832 N$27663 N$27664 "Straight Waveguide" sch_x=243 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13833 N$27665 N$27666 "Straight Waveguide" sch_x=243 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13834 N$27667 N$27668 "Straight Waveguide" sch_x=243 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13835 N$27669 N$27670 "Straight Waveguide" sch_x=243 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13836 N$27671 N$27672 "Straight Waveguide" sch_x=243 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13837 N$27673 N$27674 "Straight Waveguide" sch_x=243 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13838 N$27675 N$27676 "Straight Waveguide" sch_x=243 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13839 N$27677 N$27678 "Straight Waveguide" sch_x=243 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13840 N$27679 N$27680 "Straight Waveguide" sch_x=243 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13841 N$27681 N$27682 "Straight Waveguide" sch_x=243 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13842 N$27683 N$27684 "Straight Waveguide" sch_x=243 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13843 N$27685 N$27686 "Straight Waveguide" sch_x=243 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13844 N$27687 N$27688 "Straight Waveguide" sch_x=243 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13845 N$27689 N$27690 "Straight Waveguide" sch_x=243 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13846 N$27691 N$27692 "Straight Waveguide" sch_x=243 sch_y=-57.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13847 N$27693 N$27694 "Straight Waveguide" sch_x=241 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13848 N$27695 N$27696 "Straight Waveguide" sch_x=241 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13849 N$27697 N$27698 "Straight Waveguide" sch_x=241 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13850 N$27699 N$27700 "Straight Waveguide" sch_x=241 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13851 N$27701 N$27702 "Straight Waveguide" sch_x=241 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13852 N$27703 N$27704 "Straight Waveguide" sch_x=241 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13853 N$27705 N$27706 "Straight Waveguide" sch_x=241 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13854 N$27707 N$27708 "Straight Waveguide" sch_x=241 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13855 N$27709 N$27710 "Straight Waveguide" sch_x=241 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13856 N$27711 N$27712 "Straight Waveguide" sch_x=241 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13857 N$27713 N$27714 "Straight Waveguide" sch_x=241 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13858 N$27715 N$27716 "Straight Waveguide" sch_x=241 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13859 N$27717 N$27718 "Straight Waveguide" sch_x=241 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13860 N$27719 N$27720 "Straight Waveguide" sch_x=241 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13861 N$27721 N$27722 "Straight Waveguide" sch_x=241 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13862 N$27723 N$27724 "Straight Waveguide" sch_x=241 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13863 N$27725 N$27726 "Straight Waveguide" sch_x=241 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13864 N$27727 N$27728 "Straight Waveguide" sch_x=241 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13865 N$27729 N$27730 "Straight Waveguide" sch_x=241 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13866 N$27731 N$27732 "Straight Waveguide" sch_x=241 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13867 N$27733 N$27734 "Straight Waveguide" sch_x=241 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13868 N$27735 N$27736 "Straight Waveguide" sch_x=241 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13869 N$27737 N$27738 "Straight Waveguide" sch_x=241 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13870 N$27739 N$27740 "Straight Waveguide" sch_x=241 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13871 N$27741 N$27742 "Straight Waveguide" sch_x=241 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13872 N$27743 N$27744 "Straight Waveguide" sch_x=241 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13873 N$27745 N$27746 "Straight Waveguide" sch_x=241 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13874 N$27747 N$27748 "Straight Waveguide" sch_x=241 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13875 N$27749 N$27750 "Straight Waveguide" sch_x=241 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13876 N$27751 N$27752 "Straight Waveguide" sch_x=241 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13877 N$27753 N$27754 "Straight Waveguide" sch_x=241 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13878 N$27755 N$27756 "Straight Waveguide" sch_x=241 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13879 N$27757 N$27758 "Straight Waveguide" sch_x=241 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13880 N$27759 N$27760 "Straight Waveguide" sch_x=241 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13881 N$27761 N$27762 "Straight Waveguide" sch_x=241 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13882 N$27763 N$27764 "Straight Waveguide" sch_x=241 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13883 N$27765 N$27766 "Straight Waveguide" sch_x=241 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13884 N$27767 N$27768 "Straight Waveguide" sch_x=241 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13885 N$27769 N$27770 "Straight Waveguide" sch_x=241 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13886 N$27771 N$27772 "Straight Waveguide" sch_x=241 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13887 N$27773 N$27774 "Straight Waveguide" sch_x=241 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13888 N$27775 N$27776 "Straight Waveguide" sch_x=241 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13889 N$27777 N$27778 "Straight Waveguide" sch_x=241 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13890 N$27779 N$27780 "Straight Waveguide" sch_x=241 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13891 N$27781 N$27782 "Straight Waveguide" sch_x=241 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13892 N$27783 N$27784 "Straight Waveguide" sch_x=241 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13893 N$27785 N$27786 "Straight Waveguide" sch_x=241 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13894 N$27787 N$27788 "Straight Waveguide" sch_x=241 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13895 N$27789 N$27790 "Straight Waveguide" sch_x=241 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13896 N$27791 N$27792 "Straight Waveguide" sch_x=241 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13897 N$27793 N$27794 "Straight Waveguide" sch_x=241 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13898 N$27795 N$27796 "Straight Waveguide" sch_x=241 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13899 N$27797 N$27798 "Straight Waveguide" sch_x=241 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13900 N$27799 N$27800 "Straight Waveguide" sch_x=241 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13901 N$27801 N$27802 "Straight Waveguide" sch_x=241 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13902 N$27803 N$27804 "Straight Waveguide" sch_x=241 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13903 N$27805 N$27806 "Straight Waveguide" sch_x=241 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13904 N$27807 N$27808 "Straight Waveguide" sch_x=241 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13905 N$27809 N$27810 "Straight Waveguide" sch_x=241 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13906 N$27811 N$27812 "Straight Waveguide" sch_x=241 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13907 N$27813 N$27814 "Straight Waveguide" sch_x=241 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13908 N$27815 N$27816 "Straight Waveguide" sch_x=241 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13909 N$27817 N$27818 "Straight Waveguide" sch_x=241 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13910 N$27819 N$27820 "Straight Waveguide" sch_x=241 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13911 N$27821 N$27822 "Straight Waveguide" sch_x=241 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13912 N$27823 N$27824 "Straight Waveguide" sch_x=241 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13913 N$27825 N$27826 "Straight Waveguide" sch_x=241 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13914 N$27827 N$27828 "Straight Waveguide" sch_x=241 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13915 N$27829 N$27830 "Straight Waveguide" sch_x=241 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13916 N$27831 N$27832 "Straight Waveguide" sch_x=241 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13917 N$27833 N$27834 "Straight Waveguide" sch_x=241 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13918 N$27835 N$27836 "Straight Waveguide" sch_x=241 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13919 N$27837 N$27838 "Straight Waveguide" sch_x=241 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13920 N$27839 N$27840 "Straight Waveguide" sch_x=241 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13921 N$27841 N$27842 "Straight Waveguide" sch_x=241 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13922 N$27843 N$27844 "Straight Waveguide" sch_x=241 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13923 N$27845 N$27846 "Straight Waveguide" sch_x=241 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13924 N$27847 N$27848 "Straight Waveguide" sch_x=241 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13925 N$27849 N$27850 "Straight Waveguide" sch_x=241 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13926 N$27851 N$27852 "Straight Waveguide" sch_x=241 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13927 N$27853 N$27854 "Straight Waveguide" sch_x=241 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13928 N$27855 N$27856 "Straight Waveguide" sch_x=241 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13929 N$27857 N$27858 "Straight Waveguide" sch_x=241 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13930 N$27859 N$27860 "Straight Waveguide" sch_x=241 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13931 N$27861 N$27862 "Straight Waveguide" sch_x=241 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13932 N$27863 N$27864 "Straight Waveguide" sch_x=241 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13933 N$27865 N$27866 "Straight Waveguide" sch_x=241 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13934 N$27867 N$27868 "Straight Waveguide" sch_x=241 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13935 N$27869 N$27870 "Straight Waveguide" sch_x=241 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13936 N$27871 N$27872 "Straight Waveguide" sch_x=241 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13937 N$27873 N$27874 "Straight Waveguide" sch_x=241 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13938 N$27875 N$27876 "Straight Waveguide" sch_x=241 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13939 N$27877 N$27878 "Straight Waveguide" sch_x=241 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13940 N$27879 N$27880 "Straight Waveguide" sch_x=241 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13941 N$27881 N$27882 "Straight Waveguide" sch_x=241 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13942 N$27883 N$27884 "Straight Waveguide" sch_x=241 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13943 N$27885 N$27886 "Straight Waveguide" sch_x=241 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13944 N$27887 N$27888 "Straight Waveguide" sch_x=241 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13945 N$27889 N$27890 "Straight Waveguide" sch_x=241 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13946 N$27891 N$27892 "Straight Waveguide" sch_x=241 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13947 N$27893 N$27894 "Straight Waveguide" sch_x=241 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13948 N$27895 N$27896 "Straight Waveguide" sch_x=241 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13949 N$27897 N$27898 "Straight Waveguide" sch_x=241 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13950 N$27899 N$27900 "Straight Waveguide" sch_x=241 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13951 N$27901 N$27902 "Straight Waveguide" sch_x=241 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13952 N$27903 N$27904 "Straight Waveguide" sch_x=241 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13953 N$27905 N$27906 "Straight Waveguide" sch_x=241 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13954 N$27907 N$27908 "Straight Waveguide" sch_x=241 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13955 N$27909 N$27910 "Straight Waveguide" sch_x=241 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13956 N$27911 N$27912 "Straight Waveguide" sch_x=241 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13957 N$27913 N$27914 "Straight Waveguide" sch_x=241 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13958 N$27915 N$27916 "Straight Waveguide" sch_x=241 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13959 N$27917 N$27918 "Straight Waveguide" sch_x=241 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13960 N$27919 N$27920 "Straight Waveguide" sch_x=241 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13961 N$27921 N$27922 "Straight Waveguide" sch_x=239 sch_y=55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13962 N$27923 N$27924 "Straight Waveguide" sch_x=239 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13963 N$27925 N$27926 "Straight Waveguide" sch_x=239 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13964 N$27927 N$27928 "Straight Waveguide" sch_x=239 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13965 N$27929 N$27930 "Straight Waveguide" sch_x=239 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13966 N$27931 N$27932 "Straight Waveguide" sch_x=239 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13967 N$27933 N$27934 "Straight Waveguide" sch_x=239 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13968 N$27935 N$27936 "Straight Waveguide" sch_x=239 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13969 N$27937 N$27938 "Straight Waveguide" sch_x=239 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13970 N$27939 N$27940 "Straight Waveguide" sch_x=239 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13971 N$27941 N$27942 "Straight Waveguide" sch_x=239 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13972 N$27943 N$27944 "Straight Waveguide" sch_x=239 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13973 N$27945 N$27946 "Straight Waveguide" sch_x=239 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13974 N$27947 N$27948 "Straight Waveguide" sch_x=239 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13975 N$27949 N$27950 "Straight Waveguide" sch_x=239 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13976 N$27951 N$27952 "Straight Waveguide" sch_x=239 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13977 N$27953 N$27954 "Straight Waveguide" sch_x=239 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13978 N$27955 N$27956 "Straight Waveguide" sch_x=239 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13979 N$27957 N$27958 "Straight Waveguide" sch_x=239 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13980 N$27959 N$27960 "Straight Waveguide" sch_x=239 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13981 N$27961 N$27962 "Straight Waveguide" sch_x=239 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13982 N$27963 N$27964 "Straight Waveguide" sch_x=239 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13983 N$27965 N$27966 "Straight Waveguide" sch_x=239 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13984 N$27967 N$27968 "Straight Waveguide" sch_x=239 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13985 N$27969 N$27970 "Straight Waveguide" sch_x=239 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13986 N$27971 N$27972 "Straight Waveguide" sch_x=239 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13987 N$27973 N$27974 "Straight Waveguide" sch_x=239 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13988 N$27975 N$27976 "Straight Waveguide" sch_x=239 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13989 N$27977 N$27978 "Straight Waveguide" sch_x=239 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13990 N$27979 N$27980 "Straight Waveguide" sch_x=239 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13991 N$27981 N$27982 "Straight Waveguide" sch_x=239 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13992 N$27983 N$27984 "Straight Waveguide" sch_x=239 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13993 N$27985 N$27986 "Straight Waveguide" sch_x=239 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13994 N$27987 N$27988 "Straight Waveguide" sch_x=239 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13995 N$27989 N$27990 "Straight Waveguide" sch_x=239 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13996 N$27991 N$27992 "Straight Waveguide" sch_x=239 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13997 N$27993 N$27994 "Straight Waveguide" sch_x=239 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13998 N$27995 N$27996 "Straight Waveguide" sch_x=239 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13999 N$27997 N$27998 "Straight Waveguide" sch_x=239 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14000 N$27999 N$28000 "Straight Waveguide" sch_x=239 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14001 N$28001 N$28002 "Straight Waveguide" sch_x=239 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14002 N$28003 N$28004 "Straight Waveguide" sch_x=239 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14003 N$28005 N$28006 "Straight Waveguide" sch_x=239 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14004 N$28007 N$28008 "Straight Waveguide" sch_x=239 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14005 N$28009 N$28010 "Straight Waveguide" sch_x=239 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14006 N$28011 N$28012 "Straight Waveguide" sch_x=239 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14007 N$28013 N$28014 "Straight Waveguide" sch_x=239 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14008 N$28015 N$28016 "Straight Waveguide" sch_x=239 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14009 N$28017 N$28018 "Straight Waveguide" sch_x=239 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14010 N$28019 N$28020 "Straight Waveguide" sch_x=239 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14011 N$28021 N$28022 "Straight Waveguide" sch_x=239 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14012 N$28023 N$28024 "Straight Waveguide" sch_x=239 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14013 N$28025 N$28026 "Straight Waveguide" sch_x=239 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14014 N$28027 N$28028 "Straight Waveguide" sch_x=239 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14015 N$28029 N$28030 "Straight Waveguide" sch_x=239 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14016 N$28031 N$28032 "Straight Waveguide" sch_x=239 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14017 N$28033 N$28034 "Straight Waveguide" sch_x=239 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14018 N$28035 N$28036 "Straight Waveguide" sch_x=239 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14019 N$28037 N$28038 "Straight Waveguide" sch_x=239 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14020 N$28039 N$28040 "Straight Waveguide" sch_x=239 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14021 N$28041 N$28042 "Straight Waveguide" sch_x=239 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14022 N$28043 N$28044 "Straight Waveguide" sch_x=239 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14023 N$28045 N$28046 "Straight Waveguide" sch_x=239 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14024 N$28047 N$28048 "Straight Waveguide" sch_x=239 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14025 N$28049 N$28050 "Straight Waveguide" sch_x=239 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14026 N$28051 N$28052 "Straight Waveguide" sch_x=239 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14027 N$28053 N$28054 "Straight Waveguide" sch_x=239 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14028 N$28055 N$28056 "Straight Waveguide" sch_x=239 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14029 N$28057 N$28058 "Straight Waveguide" sch_x=239 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14030 N$28059 N$28060 "Straight Waveguide" sch_x=239 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14031 N$28061 N$28062 "Straight Waveguide" sch_x=239 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14032 N$28063 N$28064 "Straight Waveguide" sch_x=239 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14033 N$28065 N$28066 "Straight Waveguide" sch_x=239 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14034 N$28067 N$28068 "Straight Waveguide" sch_x=239 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14035 N$28069 N$28070 "Straight Waveguide" sch_x=239 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14036 N$28071 N$28072 "Straight Waveguide" sch_x=239 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14037 N$28073 N$28074 "Straight Waveguide" sch_x=239 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14038 N$28075 N$28076 "Straight Waveguide" sch_x=239 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14039 N$28077 N$28078 "Straight Waveguide" sch_x=239 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14040 N$28079 N$28080 "Straight Waveguide" sch_x=239 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14041 N$28081 N$28082 "Straight Waveguide" sch_x=239 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14042 N$28083 N$28084 "Straight Waveguide" sch_x=239 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14043 N$28085 N$28086 "Straight Waveguide" sch_x=239 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14044 N$28087 N$28088 "Straight Waveguide" sch_x=239 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14045 N$28089 N$28090 "Straight Waveguide" sch_x=239 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14046 N$28091 N$28092 "Straight Waveguide" sch_x=239 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14047 N$28093 N$28094 "Straight Waveguide" sch_x=239 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14048 N$28095 N$28096 "Straight Waveguide" sch_x=239 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14049 N$28097 N$28098 "Straight Waveguide" sch_x=239 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14050 N$28099 N$28100 "Straight Waveguide" sch_x=239 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14051 N$28101 N$28102 "Straight Waveguide" sch_x=239 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14052 N$28103 N$28104 "Straight Waveguide" sch_x=239 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14053 N$28105 N$28106 "Straight Waveguide" sch_x=239 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14054 N$28107 N$28108 "Straight Waveguide" sch_x=239 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14055 N$28109 N$28110 "Straight Waveguide" sch_x=239 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14056 N$28111 N$28112 "Straight Waveguide" sch_x=239 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14057 N$28113 N$28114 "Straight Waveguide" sch_x=239 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14058 N$28115 N$28116 "Straight Waveguide" sch_x=239 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14059 N$28117 N$28118 "Straight Waveguide" sch_x=239 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14060 N$28119 N$28120 "Straight Waveguide" sch_x=239 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14061 N$28121 N$28122 "Straight Waveguide" sch_x=239 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14062 N$28123 N$28124 "Straight Waveguide" sch_x=239 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14063 N$28125 N$28126 "Straight Waveguide" sch_x=239 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14064 N$28127 N$28128 "Straight Waveguide" sch_x=239 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14065 N$28129 N$28130 "Straight Waveguide" sch_x=239 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14066 N$28131 N$28132 "Straight Waveguide" sch_x=239 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14067 N$28133 N$28134 "Straight Waveguide" sch_x=239 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14068 N$28135 N$28136 "Straight Waveguide" sch_x=239 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14069 N$28137 N$28138 "Straight Waveguide" sch_x=239 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14070 N$28139 N$28140 "Straight Waveguide" sch_x=239 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14071 N$28141 N$28142 "Straight Waveguide" sch_x=239 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14072 N$28143 N$28144 "Straight Waveguide" sch_x=239 sch_y=-55.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14073 N$28145 N$28146 "Straight Waveguide" sch_x=237 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14074 N$28147 N$28148 "Straight Waveguide" sch_x=237 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14075 N$28149 N$28150 "Straight Waveguide" sch_x=237 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14076 N$28151 N$28152 "Straight Waveguide" sch_x=237 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14077 N$28153 N$28154 "Straight Waveguide" sch_x=237 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14078 N$28155 N$28156 "Straight Waveguide" sch_x=237 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14079 N$28157 N$28158 "Straight Waveguide" sch_x=237 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14080 N$28159 N$28160 "Straight Waveguide" sch_x=237 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14081 N$28161 N$28162 "Straight Waveguide" sch_x=237 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14082 N$28163 N$28164 "Straight Waveguide" sch_x=237 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14083 N$28165 N$28166 "Straight Waveguide" sch_x=237 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14084 N$28167 N$28168 "Straight Waveguide" sch_x=237 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14085 N$28169 N$28170 "Straight Waveguide" sch_x=237 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14086 N$28171 N$28172 "Straight Waveguide" sch_x=237 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14087 N$28173 N$28174 "Straight Waveguide" sch_x=237 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14088 N$28175 N$28176 "Straight Waveguide" sch_x=237 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14089 N$28177 N$28178 "Straight Waveguide" sch_x=237 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14090 N$28179 N$28180 "Straight Waveguide" sch_x=237 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14091 N$28181 N$28182 "Straight Waveguide" sch_x=237 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14092 N$28183 N$28184 "Straight Waveguide" sch_x=237 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14093 N$28185 N$28186 "Straight Waveguide" sch_x=237 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14094 N$28187 N$28188 "Straight Waveguide" sch_x=237 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14095 N$28189 N$28190 "Straight Waveguide" sch_x=237 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14096 N$28191 N$28192 "Straight Waveguide" sch_x=237 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14097 N$28193 N$28194 "Straight Waveguide" sch_x=237 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14098 N$28195 N$28196 "Straight Waveguide" sch_x=237 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14099 N$28197 N$28198 "Straight Waveguide" sch_x=237 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14100 N$28199 N$28200 "Straight Waveguide" sch_x=237 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14101 N$28201 N$28202 "Straight Waveguide" sch_x=237 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14102 N$28203 N$28204 "Straight Waveguide" sch_x=237 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14103 N$28205 N$28206 "Straight Waveguide" sch_x=237 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14104 N$28207 N$28208 "Straight Waveguide" sch_x=237 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14105 N$28209 N$28210 "Straight Waveguide" sch_x=237 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14106 N$28211 N$28212 "Straight Waveguide" sch_x=237 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14107 N$28213 N$28214 "Straight Waveguide" sch_x=237 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14108 N$28215 N$28216 "Straight Waveguide" sch_x=237 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14109 N$28217 N$28218 "Straight Waveguide" sch_x=237 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14110 N$28219 N$28220 "Straight Waveguide" sch_x=237 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14111 N$28221 N$28222 "Straight Waveguide" sch_x=237 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14112 N$28223 N$28224 "Straight Waveguide" sch_x=237 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14113 N$28225 N$28226 "Straight Waveguide" sch_x=237 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14114 N$28227 N$28228 "Straight Waveguide" sch_x=237 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14115 N$28229 N$28230 "Straight Waveguide" sch_x=237 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14116 N$28231 N$28232 "Straight Waveguide" sch_x=237 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14117 N$28233 N$28234 "Straight Waveguide" sch_x=237 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14118 N$28235 N$28236 "Straight Waveguide" sch_x=237 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14119 N$28237 N$28238 "Straight Waveguide" sch_x=237 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14120 N$28239 N$28240 "Straight Waveguide" sch_x=237 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14121 N$28241 N$28242 "Straight Waveguide" sch_x=237 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14122 N$28243 N$28244 "Straight Waveguide" sch_x=237 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14123 N$28245 N$28246 "Straight Waveguide" sch_x=237 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14124 N$28247 N$28248 "Straight Waveguide" sch_x=237 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14125 N$28249 N$28250 "Straight Waveguide" sch_x=237 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14126 N$28251 N$28252 "Straight Waveguide" sch_x=237 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14127 N$28253 N$28254 "Straight Waveguide" sch_x=237 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14128 N$28255 N$28256 "Straight Waveguide" sch_x=237 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14129 N$28257 N$28258 "Straight Waveguide" sch_x=237 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14130 N$28259 N$28260 "Straight Waveguide" sch_x=237 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14131 N$28261 N$28262 "Straight Waveguide" sch_x=237 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14132 N$28263 N$28264 "Straight Waveguide" sch_x=237 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14133 N$28265 N$28266 "Straight Waveguide" sch_x=237 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14134 N$28267 N$28268 "Straight Waveguide" sch_x=237 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14135 N$28269 N$28270 "Straight Waveguide" sch_x=237 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14136 N$28271 N$28272 "Straight Waveguide" sch_x=237 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14137 N$28273 N$28274 "Straight Waveguide" sch_x=237 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14138 N$28275 N$28276 "Straight Waveguide" sch_x=237 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14139 N$28277 N$28278 "Straight Waveguide" sch_x=237 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14140 N$28279 N$28280 "Straight Waveguide" sch_x=237 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14141 N$28281 N$28282 "Straight Waveguide" sch_x=237 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14142 N$28283 N$28284 "Straight Waveguide" sch_x=237 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14143 N$28285 N$28286 "Straight Waveguide" sch_x=237 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14144 N$28287 N$28288 "Straight Waveguide" sch_x=237 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14145 N$28289 N$28290 "Straight Waveguide" sch_x=237 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14146 N$28291 N$28292 "Straight Waveguide" sch_x=237 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14147 N$28293 N$28294 "Straight Waveguide" sch_x=237 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14148 N$28295 N$28296 "Straight Waveguide" sch_x=237 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14149 N$28297 N$28298 "Straight Waveguide" sch_x=237 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14150 N$28299 N$28300 "Straight Waveguide" sch_x=237 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14151 N$28301 N$28302 "Straight Waveguide" sch_x=237 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14152 N$28303 N$28304 "Straight Waveguide" sch_x=237 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14153 N$28305 N$28306 "Straight Waveguide" sch_x=237 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14154 N$28307 N$28308 "Straight Waveguide" sch_x=237 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14155 N$28309 N$28310 "Straight Waveguide" sch_x=237 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14156 N$28311 N$28312 "Straight Waveguide" sch_x=237 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14157 N$28313 N$28314 "Straight Waveguide" sch_x=237 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14158 N$28315 N$28316 "Straight Waveguide" sch_x=237 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14159 N$28317 N$28318 "Straight Waveguide" sch_x=237 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14160 N$28319 N$28320 "Straight Waveguide" sch_x=237 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14161 N$28321 N$28322 "Straight Waveguide" sch_x=237 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14162 N$28323 N$28324 "Straight Waveguide" sch_x=237 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14163 N$28325 N$28326 "Straight Waveguide" sch_x=237 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14164 N$28327 N$28328 "Straight Waveguide" sch_x=237 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14165 N$28329 N$28330 "Straight Waveguide" sch_x=237 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14166 N$28331 N$28332 "Straight Waveguide" sch_x=237 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14167 N$28333 N$28334 "Straight Waveguide" sch_x=237 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14168 N$28335 N$28336 "Straight Waveguide" sch_x=237 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14169 N$28337 N$28338 "Straight Waveguide" sch_x=237 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14170 N$28339 N$28340 "Straight Waveguide" sch_x=237 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14171 N$28341 N$28342 "Straight Waveguide" sch_x=237 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14172 N$28343 N$28344 "Straight Waveguide" sch_x=237 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14173 N$28345 N$28346 "Straight Waveguide" sch_x=237 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14174 N$28347 N$28348 "Straight Waveguide" sch_x=237 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14175 N$28349 N$28350 "Straight Waveguide" sch_x=237 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14176 N$28351 N$28352 "Straight Waveguide" sch_x=237 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14177 N$28353 N$28354 "Straight Waveguide" sch_x=237 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14178 N$28355 N$28356 "Straight Waveguide" sch_x=237 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14179 N$28357 N$28358 "Straight Waveguide" sch_x=237 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14180 N$28359 N$28360 "Straight Waveguide" sch_x=237 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14181 N$28361 N$28362 "Straight Waveguide" sch_x=237 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14182 N$28363 N$28364 "Straight Waveguide" sch_x=237 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14183 N$28365 N$28366 "Straight Waveguide" sch_x=235 sch_y=53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14184 N$28367 N$28368 "Straight Waveguide" sch_x=235 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14185 N$28369 N$28370 "Straight Waveguide" sch_x=235 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14186 N$28371 N$28372 "Straight Waveguide" sch_x=235 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14187 N$28373 N$28374 "Straight Waveguide" sch_x=235 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14188 N$28375 N$28376 "Straight Waveguide" sch_x=235 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14189 N$28377 N$28378 "Straight Waveguide" sch_x=235 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14190 N$28379 N$28380 "Straight Waveguide" sch_x=235 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14191 N$28381 N$28382 "Straight Waveguide" sch_x=235 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14192 N$28383 N$28384 "Straight Waveguide" sch_x=235 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14193 N$28385 N$28386 "Straight Waveguide" sch_x=235 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14194 N$28387 N$28388 "Straight Waveguide" sch_x=235 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14195 N$28389 N$28390 "Straight Waveguide" sch_x=235 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14196 N$28391 N$28392 "Straight Waveguide" sch_x=235 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14197 N$28393 N$28394 "Straight Waveguide" sch_x=235 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14198 N$28395 N$28396 "Straight Waveguide" sch_x=235 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14199 N$28397 N$28398 "Straight Waveguide" sch_x=235 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14200 N$28399 N$28400 "Straight Waveguide" sch_x=235 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14201 N$28401 N$28402 "Straight Waveguide" sch_x=235 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14202 N$28403 N$28404 "Straight Waveguide" sch_x=235 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14203 N$28405 N$28406 "Straight Waveguide" sch_x=235 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14204 N$28407 N$28408 "Straight Waveguide" sch_x=235 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14205 N$28409 N$28410 "Straight Waveguide" sch_x=235 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14206 N$28411 N$28412 "Straight Waveguide" sch_x=235 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14207 N$28413 N$28414 "Straight Waveguide" sch_x=235 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14208 N$28415 N$28416 "Straight Waveguide" sch_x=235 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14209 N$28417 N$28418 "Straight Waveguide" sch_x=235 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14210 N$28419 N$28420 "Straight Waveguide" sch_x=235 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14211 N$28421 N$28422 "Straight Waveguide" sch_x=235 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14212 N$28423 N$28424 "Straight Waveguide" sch_x=235 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14213 N$28425 N$28426 "Straight Waveguide" sch_x=235 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14214 N$28427 N$28428 "Straight Waveguide" sch_x=235 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14215 N$28429 N$28430 "Straight Waveguide" sch_x=235 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14216 N$28431 N$28432 "Straight Waveguide" sch_x=235 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14217 N$28433 N$28434 "Straight Waveguide" sch_x=235 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14218 N$28435 N$28436 "Straight Waveguide" sch_x=235 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14219 N$28437 N$28438 "Straight Waveguide" sch_x=235 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14220 N$28439 N$28440 "Straight Waveguide" sch_x=235 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14221 N$28441 N$28442 "Straight Waveguide" sch_x=235 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14222 N$28443 N$28444 "Straight Waveguide" sch_x=235 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14223 N$28445 N$28446 "Straight Waveguide" sch_x=235 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14224 N$28447 N$28448 "Straight Waveguide" sch_x=235 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14225 N$28449 N$28450 "Straight Waveguide" sch_x=235 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14226 N$28451 N$28452 "Straight Waveguide" sch_x=235 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14227 N$28453 N$28454 "Straight Waveguide" sch_x=235 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14228 N$28455 N$28456 "Straight Waveguide" sch_x=235 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14229 N$28457 N$28458 "Straight Waveguide" sch_x=235 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14230 N$28459 N$28460 "Straight Waveguide" sch_x=235 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14231 N$28461 N$28462 "Straight Waveguide" sch_x=235 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14232 N$28463 N$28464 "Straight Waveguide" sch_x=235 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14233 N$28465 N$28466 "Straight Waveguide" sch_x=235 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14234 N$28467 N$28468 "Straight Waveguide" sch_x=235 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14235 N$28469 N$28470 "Straight Waveguide" sch_x=235 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14236 N$28471 N$28472 "Straight Waveguide" sch_x=235 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14237 N$28473 N$28474 "Straight Waveguide" sch_x=235 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14238 N$28475 N$28476 "Straight Waveguide" sch_x=235 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14239 N$28477 N$28478 "Straight Waveguide" sch_x=235 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14240 N$28479 N$28480 "Straight Waveguide" sch_x=235 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14241 N$28481 N$28482 "Straight Waveguide" sch_x=235 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14242 N$28483 N$28484 "Straight Waveguide" sch_x=235 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14243 N$28485 N$28486 "Straight Waveguide" sch_x=235 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14244 N$28487 N$28488 "Straight Waveguide" sch_x=235 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14245 N$28489 N$28490 "Straight Waveguide" sch_x=235 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14246 N$28491 N$28492 "Straight Waveguide" sch_x=235 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14247 N$28493 N$28494 "Straight Waveguide" sch_x=235 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14248 N$28495 N$28496 "Straight Waveguide" sch_x=235 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14249 N$28497 N$28498 "Straight Waveguide" sch_x=235 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14250 N$28499 N$28500 "Straight Waveguide" sch_x=235 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14251 N$28501 N$28502 "Straight Waveguide" sch_x=235 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14252 N$28503 N$28504 "Straight Waveguide" sch_x=235 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14253 N$28505 N$28506 "Straight Waveguide" sch_x=235 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14254 N$28507 N$28508 "Straight Waveguide" sch_x=235 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14255 N$28509 N$28510 "Straight Waveguide" sch_x=235 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14256 N$28511 N$28512 "Straight Waveguide" sch_x=235 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14257 N$28513 N$28514 "Straight Waveguide" sch_x=235 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14258 N$28515 N$28516 "Straight Waveguide" sch_x=235 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14259 N$28517 N$28518 "Straight Waveguide" sch_x=235 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14260 N$28519 N$28520 "Straight Waveguide" sch_x=235 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14261 N$28521 N$28522 "Straight Waveguide" sch_x=235 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14262 N$28523 N$28524 "Straight Waveguide" sch_x=235 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14263 N$28525 N$28526 "Straight Waveguide" sch_x=235 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14264 N$28527 N$28528 "Straight Waveguide" sch_x=235 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14265 N$28529 N$28530 "Straight Waveguide" sch_x=235 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14266 N$28531 N$28532 "Straight Waveguide" sch_x=235 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14267 N$28533 N$28534 "Straight Waveguide" sch_x=235 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14268 N$28535 N$28536 "Straight Waveguide" sch_x=235 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14269 N$28537 N$28538 "Straight Waveguide" sch_x=235 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14270 N$28539 N$28540 "Straight Waveguide" sch_x=235 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14271 N$28541 N$28542 "Straight Waveguide" sch_x=235 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14272 N$28543 N$28544 "Straight Waveguide" sch_x=235 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14273 N$28545 N$28546 "Straight Waveguide" sch_x=235 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14274 N$28547 N$28548 "Straight Waveguide" sch_x=235 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14275 N$28549 N$28550 "Straight Waveguide" sch_x=235 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14276 N$28551 N$28552 "Straight Waveguide" sch_x=235 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14277 N$28553 N$28554 "Straight Waveguide" sch_x=235 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14278 N$28555 N$28556 "Straight Waveguide" sch_x=235 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14279 N$28557 N$28558 "Straight Waveguide" sch_x=235 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14280 N$28559 N$28560 "Straight Waveguide" sch_x=235 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14281 N$28561 N$28562 "Straight Waveguide" sch_x=235 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14282 N$28563 N$28564 "Straight Waveguide" sch_x=235 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14283 N$28565 N$28566 "Straight Waveguide" sch_x=235 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14284 N$28567 N$28568 "Straight Waveguide" sch_x=235 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14285 N$28569 N$28570 "Straight Waveguide" sch_x=235 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14286 N$28571 N$28572 "Straight Waveguide" sch_x=235 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14287 N$28573 N$28574 "Straight Waveguide" sch_x=235 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14288 N$28575 N$28576 "Straight Waveguide" sch_x=235 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14289 N$28577 N$28578 "Straight Waveguide" sch_x=235 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14290 N$28579 N$28580 "Straight Waveguide" sch_x=235 sch_y=-53.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14291 N$28581 N$28582 "Straight Waveguide" sch_x=233 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14292 N$28583 N$28584 "Straight Waveguide" sch_x=233 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14293 N$28585 N$28586 "Straight Waveguide" sch_x=233 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14294 N$28587 N$28588 "Straight Waveguide" sch_x=233 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14295 N$28589 N$28590 "Straight Waveguide" sch_x=233 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14296 N$28591 N$28592 "Straight Waveguide" sch_x=233 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14297 N$28593 N$28594 "Straight Waveguide" sch_x=233 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14298 N$28595 N$28596 "Straight Waveguide" sch_x=233 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14299 N$28597 N$28598 "Straight Waveguide" sch_x=233 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14300 N$28599 N$28600 "Straight Waveguide" sch_x=233 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14301 N$28601 N$28602 "Straight Waveguide" sch_x=233 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14302 N$28603 N$28604 "Straight Waveguide" sch_x=233 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14303 N$28605 N$28606 "Straight Waveguide" sch_x=233 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14304 N$28607 N$28608 "Straight Waveguide" sch_x=233 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14305 N$28609 N$28610 "Straight Waveguide" sch_x=233 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14306 N$28611 N$28612 "Straight Waveguide" sch_x=233 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14307 N$28613 N$28614 "Straight Waveguide" sch_x=233 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14308 N$28615 N$28616 "Straight Waveguide" sch_x=233 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14309 N$28617 N$28618 "Straight Waveguide" sch_x=233 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14310 N$28619 N$28620 "Straight Waveguide" sch_x=233 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14311 N$28621 N$28622 "Straight Waveguide" sch_x=233 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14312 N$28623 N$28624 "Straight Waveguide" sch_x=233 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14313 N$28625 N$28626 "Straight Waveguide" sch_x=233 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14314 N$28627 N$28628 "Straight Waveguide" sch_x=233 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14315 N$28629 N$28630 "Straight Waveguide" sch_x=233 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14316 N$28631 N$28632 "Straight Waveguide" sch_x=233 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14317 N$28633 N$28634 "Straight Waveguide" sch_x=233 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14318 N$28635 N$28636 "Straight Waveguide" sch_x=233 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14319 N$28637 N$28638 "Straight Waveguide" sch_x=233 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14320 N$28639 N$28640 "Straight Waveguide" sch_x=233 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14321 N$28641 N$28642 "Straight Waveguide" sch_x=233 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14322 N$28643 N$28644 "Straight Waveguide" sch_x=233 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14323 N$28645 N$28646 "Straight Waveguide" sch_x=233 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14324 N$28647 N$28648 "Straight Waveguide" sch_x=233 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14325 N$28649 N$28650 "Straight Waveguide" sch_x=233 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14326 N$28651 N$28652 "Straight Waveguide" sch_x=233 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14327 N$28653 N$28654 "Straight Waveguide" sch_x=233 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14328 N$28655 N$28656 "Straight Waveguide" sch_x=233 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14329 N$28657 N$28658 "Straight Waveguide" sch_x=233 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14330 N$28659 N$28660 "Straight Waveguide" sch_x=233 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14331 N$28661 N$28662 "Straight Waveguide" sch_x=233 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14332 N$28663 N$28664 "Straight Waveguide" sch_x=233 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14333 N$28665 N$28666 "Straight Waveguide" sch_x=233 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14334 N$28667 N$28668 "Straight Waveguide" sch_x=233 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14335 N$28669 N$28670 "Straight Waveguide" sch_x=233 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14336 N$28671 N$28672 "Straight Waveguide" sch_x=233 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14337 N$28673 N$28674 "Straight Waveguide" sch_x=233 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14338 N$28675 N$28676 "Straight Waveguide" sch_x=233 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14339 N$28677 N$28678 "Straight Waveguide" sch_x=233 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14340 N$28679 N$28680 "Straight Waveguide" sch_x=233 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14341 N$28681 N$28682 "Straight Waveguide" sch_x=233 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14342 N$28683 N$28684 "Straight Waveguide" sch_x=233 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14343 N$28685 N$28686 "Straight Waveguide" sch_x=233 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14344 N$28687 N$28688 "Straight Waveguide" sch_x=233 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14345 N$28689 N$28690 "Straight Waveguide" sch_x=233 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14346 N$28691 N$28692 "Straight Waveguide" sch_x=233 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14347 N$28693 N$28694 "Straight Waveguide" sch_x=233 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14348 N$28695 N$28696 "Straight Waveguide" sch_x=233 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14349 N$28697 N$28698 "Straight Waveguide" sch_x=233 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14350 N$28699 N$28700 "Straight Waveguide" sch_x=233 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14351 N$28701 N$28702 "Straight Waveguide" sch_x=233 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14352 N$28703 N$28704 "Straight Waveguide" sch_x=233 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14353 N$28705 N$28706 "Straight Waveguide" sch_x=233 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14354 N$28707 N$28708 "Straight Waveguide" sch_x=233 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14355 N$28709 N$28710 "Straight Waveguide" sch_x=233 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14356 N$28711 N$28712 "Straight Waveguide" sch_x=233 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14357 N$28713 N$28714 "Straight Waveguide" sch_x=233 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14358 N$28715 N$28716 "Straight Waveguide" sch_x=233 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14359 N$28717 N$28718 "Straight Waveguide" sch_x=233 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14360 N$28719 N$28720 "Straight Waveguide" sch_x=233 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14361 N$28721 N$28722 "Straight Waveguide" sch_x=233 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14362 N$28723 N$28724 "Straight Waveguide" sch_x=233 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14363 N$28725 N$28726 "Straight Waveguide" sch_x=233 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14364 N$28727 N$28728 "Straight Waveguide" sch_x=233 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14365 N$28729 N$28730 "Straight Waveguide" sch_x=233 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14366 N$28731 N$28732 "Straight Waveguide" sch_x=233 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14367 N$28733 N$28734 "Straight Waveguide" sch_x=233 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14368 N$28735 N$28736 "Straight Waveguide" sch_x=233 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14369 N$28737 N$28738 "Straight Waveguide" sch_x=233 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14370 N$28739 N$28740 "Straight Waveguide" sch_x=233 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14371 N$28741 N$28742 "Straight Waveguide" sch_x=233 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14372 N$28743 N$28744 "Straight Waveguide" sch_x=233 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14373 N$28745 N$28746 "Straight Waveguide" sch_x=233 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14374 N$28747 N$28748 "Straight Waveguide" sch_x=233 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14375 N$28749 N$28750 "Straight Waveguide" sch_x=233 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14376 N$28751 N$28752 "Straight Waveguide" sch_x=233 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14377 N$28753 N$28754 "Straight Waveguide" sch_x=233 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14378 N$28755 N$28756 "Straight Waveguide" sch_x=233 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14379 N$28757 N$28758 "Straight Waveguide" sch_x=233 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14380 N$28759 N$28760 "Straight Waveguide" sch_x=233 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14381 N$28761 N$28762 "Straight Waveguide" sch_x=233 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14382 N$28763 N$28764 "Straight Waveguide" sch_x=233 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14383 N$28765 N$28766 "Straight Waveguide" sch_x=233 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14384 N$28767 N$28768 "Straight Waveguide" sch_x=233 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14385 N$28769 N$28770 "Straight Waveguide" sch_x=233 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14386 N$28771 N$28772 "Straight Waveguide" sch_x=233 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14387 N$28773 N$28774 "Straight Waveguide" sch_x=233 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14388 N$28775 N$28776 "Straight Waveguide" sch_x=233 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14389 N$28777 N$28778 "Straight Waveguide" sch_x=233 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14390 N$28779 N$28780 "Straight Waveguide" sch_x=233 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14391 N$28781 N$28782 "Straight Waveguide" sch_x=233 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14392 N$28783 N$28784 "Straight Waveguide" sch_x=233 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14393 N$28785 N$28786 "Straight Waveguide" sch_x=233 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14394 N$28787 N$28788 "Straight Waveguide" sch_x=233 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14395 N$28789 N$28790 "Straight Waveguide" sch_x=233 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14396 N$28791 N$28792 "Straight Waveguide" sch_x=233 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14397 N$28793 N$28794 "Straight Waveguide" sch_x=231 sch_y=51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14398 N$28795 N$28796 "Straight Waveguide" sch_x=231 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14399 N$28797 N$28798 "Straight Waveguide" sch_x=231 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14400 N$28799 N$28800 "Straight Waveguide" sch_x=231 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14401 N$28801 N$28802 "Straight Waveguide" sch_x=231 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14402 N$28803 N$28804 "Straight Waveguide" sch_x=231 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14403 N$28805 N$28806 "Straight Waveguide" sch_x=231 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14404 N$28807 N$28808 "Straight Waveguide" sch_x=231 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14405 N$28809 N$28810 "Straight Waveguide" sch_x=231 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14406 N$28811 N$28812 "Straight Waveguide" sch_x=231 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14407 N$28813 N$28814 "Straight Waveguide" sch_x=231 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14408 N$28815 N$28816 "Straight Waveguide" sch_x=231 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14409 N$28817 N$28818 "Straight Waveguide" sch_x=231 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14410 N$28819 N$28820 "Straight Waveguide" sch_x=231 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14411 N$28821 N$28822 "Straight Waveguide" sch_x=231 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14412 N$28823 N$28824 "Straight Waveguide" sch_x=231 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14413 N$28825 N$28826 "Straight Waveguide" sch_x=231 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14414 N$28827 N$28828 "Straight Waveguide" sch_x=231 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14415 N$28829 N$28830 "Straight Waveguide" sch_x=231 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14416 N$28831 N$28832 "Straight Waveguide" sch_x=231 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14417 N$28833 N$28834 "Straight Waveguide" sch_x=231 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14418 N$28835 N$28836 "Straight Waveguide" sch_x=231 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14419 N$28837 N$28838 "Straight Waveguide" sch_x=231 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14420 N$28839 N$28840 "Straight Waveguide" sch_x=231 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14421 N$28841 N$28842 "Straight Waveguide" sch_x=231 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14422 N$28843 N$28844 "Straight Waveguide" sch_x=231 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14423 N$28845 N$28846 "Straight Waveguide" sch_x=231 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14424 N$28847 N$28848 "Straight Waveguide" sch_x=231 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14425 N$28849 N$28850 "Straight Waveguide" sch_x=231 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14426 N$28851 N$28852 "Straight Waveguide" sch_x=231 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14427 N$28853 N$28854 "Straight Waveguide" sch_x=231 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14428 N$28855 N$28856 "Straight Waveguide" sch_x=231 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14429 N$28857 N$28858 "Straight Waveguide" sch_x=231 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14430 N$28859 N$28860 "Straight Waveguide" sch_x=231 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14431 N$28861 N$28862 "Straight Waveguide" sch_x=231 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14432 N$28863 N$28864 "Straight Waveguide" sch_x=231 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14433 N$28865 N$28866 "Straight Waveguide" sch_x=231 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14434 N$28867 N$28868 "Straight Waveguide" sch_x=231 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14435 N$28869 N$28870 "Straight Waveguide" sch_x=231 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14436 N$28871 N$28872 "Straight Waveguide" sch_x=231 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14437 N$28873 N$28874 "Straight Waveguide" sch_x=231 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14438 N$28875 N$28876 "Straight Waveguide" sch_x=231 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14439 N$28877 N$28878 "Straight Waveguide" sch_x=231 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14440 N$28879 N$28880 "Straight Waveguide" sch_x=231 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14441 N$28881 N$28882 "Straight Waveguide" sch_x=231 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14442 N$28883 N$28884 "Straight Waveguide" sch_x=231 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14443 N$28885 N$28886 "Straight Waveguide" sch_x=231 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14444 N$28887 N$28888 "Straight Waveguide" sch_x=231 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14445 N$28889 N$28890 "Straight Waveguide" sch_x=231 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14446 N$28891 N$28892 "Straight Waveguide" sch_x=231 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14447 N$28893 N$28894 "Straight Waveguide" sch_x=231 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14448 N$28895 N$28896 "Straight Waveguide" sch_x=231 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14449 N$28897 N$28898 "Straight Waveguide" sch_x=231 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14450 N$28899 N$28900 "Straight Waveguide" sch_x=231 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14451 N$28901 N$28902 "Straight Waveguide" sch_x=231 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14452 N$28903 N$28904 "Straight Waveguide" sch_x=231 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14453 N$28905 N$28906 "Straight Waveguide" sch_x=231 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14454 N$28907 N$28908 "Straight Waveguide" sch_x=231 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14455 N$28909 N$28910 "Straight Waveguide" sch_x=231 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14456 N$28911 N$28912 "Straight Waveguide" sch_x=231 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14457 N$28913 N$28914 "Straight Waveguide" sch_x=231 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14458 N$28915 N$28916 "Straight Waveguide" sch_x=231 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14459 N$28917 N$28918 "Straight Waveguide" sch_x=231 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14460 N$28919 N$28920 "Straight Waveguide" sch_x=231 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14461 N$28921 N$28922 "Straight Waveguide" sch_x=231 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14462 N$28923 N$28924 "Straight Waveguide" sch_x=231 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14463 N$28925 N$28926 "Straight Waveguide" sch_x=231 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14464 N$28927 N$28928 "Straight Waveguide" sch_x=231 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14465 N$28929 N$28930 "Straight Waveguide" sch_x=231 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14466 N$28931 N$28932 "Straight Waveguide" sch_x=231 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14467 N$28933 N$28934 "Straight Waveguide" sch_x=231 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14468 N$28935 N$28936 "Straight Waveguide" sch_x=231 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14469 N$28937 N$28938 "Straight Waveguide" sch_x=231 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14470 N$28939 N$28940 "Straight Waveguide" sch_x=231 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14471 N$28941 N$28942 "Straight Waveguide" sch_x=231 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14472 N$28943 N$28944 "Straight Waveguide" sch_x=231 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14473 N$28945 N$28946 "Straight Waveguide" sch_x=231 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14474 N$28947 N$28948 "Straight Waveguide" sch_x=231 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14475 N$28949 N$28950 "Straight Waveguide" sch_x=231 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14476 N$28951 N$28952 "Straight Waveguide" sch_x=231 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14477 N$28953 N$28954 "Straight Waveguide" sch_x=231 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14478 N$28955 N$28956 "Straight Waveguide" sch_x=231 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14479 N$28957 N$28958 "Straight Waveguide" sch_x=231 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14480 N$28959 N$28960 "Straight Waveguide" sch_x=231 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14481 N$28961 N$28962 "Straight Waveguide" sch_x=231 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14482 N$28963 N$28964 "Straight Waveguide" sch_x=231 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14483 N$28965 N$28966 "Straight Waveguide" sch_x=231 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14484 N$28967 N$28968 "Straight Waveguide" sch_x=231 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14485 N$28969 N$28970 "Straight Waveguide" sch_x=231 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14486 N$28971 N$28972 "Straight Waveguide" sch_x=231 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14487 N$28973 N$28974 "Straight Waveguide" sch_x=231 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14488 N$28975 N$28976 "Straight Waveguide" sch_x=231 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14489 N$28977 N$28978 "Straight Waveguide" sch_x=231 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14490 N$28979 N$28980 "Straight Waveguide" sch_x=231 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14491 N$28981 N$28982 "Straight Waveguide" sch_x=231 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14492 N$28983 N$28984 "Straight Waveguide" sch_x=231 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14493 N$28985 N$28986 "Straight Waveguide" sch_x=231 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14494 N$28987 N$28988 "Straight Waveguide" sch_x=231 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14495 N$28989 N$28990 "Straight Waveguide" sch_x=231 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14496 N$28991 N$28992 "Straight Waveguide" sch_x=231 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14497 N$28993 N$28994 "Straight Waveguide" sch_x=231 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14498 N$28995 N$28996 "Straight Waveguide" sch_x=231 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14499 N$28997 N$28998 "Straight Waveguide" sch_x=231 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14500 N$28999 N$29000 "Straight Waveguide" sch_x=231 sch_y=-51.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14501 N$29001 N$29002 "Straight Waveguide" sch_x=229 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14502 N$29003 N$29004 "Straight Waveguide" sch_x=229 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14503 N$29005 N$29006 "Straight Waveguide" sch_x=229 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14504 N$29007 N$29008 "Straight Waveguide" sch_x=229 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14505 N$29009 N$29010 "Straight Waveguide" sch_x=229 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14506 N$29011 N$29012 "Straight Waveguide" sch_x=229 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14507 N$29013 N$29014 "Straight Waveguide" sch_x=229 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14508 N$29015 N$29016 "Straight Waveguide" sch_x=229 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14509 N$29017 N$29018 "Straight Waveguide" sch_x=229 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14510 N$29019 N$29020 "Straight Waveguide" sch_x=229 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14511 N$29021 N$29022 "Straight Waveguide" sch_x=229 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14512 N$29023 N$29024 "Straight Waveguide" sch_x=229 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14513 N$29025 N$29026 "Straight Waveguide" sch_x=229 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14514 N$29027 N$29028 "Straight Waveguide" sch_x=229 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14515 N$29029 N$29030 "Straight Waveguide" sch_x=229 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14516 N$29031 N$29032 "Straight Waveguide" sch_x=229 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14517 N$29033 N$29034 "Straight Waveguide" sch_x=229 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14518 N$29035 N$29036 "Straight Waveguide" sch_x=229 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14519 N$29037 N$29038 "Straight Waveguide" sch_x=229 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14520 N$29039 N$29040 "Straight Waveguide" sch_x=229 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14521 N$29041 N$29042 "Straight Waveguide" sch_x=229 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14522 N$29043 N$29044 "Straight Waveguide" sch_x=229 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14523 N$29045 N$29046 "Straight Waveguide" sch_x=229 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14524 N$29047 N$29048 "Straight Waveguide" sch_x=229 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14525 N$29049 N$29050 "Straight Waveguide" sch_x=229 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14526 N$29051 N$29052 "Straight Waveguide" sch_x=229 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14527 N$29053 N$29054 "Straight Waveguide" sch_x=229 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14528 N$29055 N$29056 "Straight Waveguide" sch_x=229 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14529 N$29057 N$29058 "Straight Waveguide" sch_x=229 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14530 N$29059 N$29060 "Straight Waveguide" sch_x=229 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14531 N$29061 N$29062 "Straight Waveguide" sch_x=229 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14532 N$29063 N$29064 "Straight Waveguide" sch_x=229 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14533 N$29065 N$29066 "Straight Waveguide" sch_x=229 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14534 N$29067 N$29068 "Straight Waveguide" sch_x=229 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14535 N$29069 N$29070 "Straight Waveguide" sch_x=229 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14536 N$29071 N$29072 "Straight Waveguide" sch_x=229 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14537 N$29073 N$29074 "Straight Waveguide" sch_x=229 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14538 N$29075 N$29076 "Straight Waveguide" sch_x=229 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14539 N$29077 N$29078 "Straight Waveguide" sch_x=229 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14540 N$29079 N$29080 "Straight Waveguide" sch_x=229 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14541 N$29081 N$29082 "Straight Waveguide" sch_x=229 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14542 N$29083 N$29084 "Straight Waveguide" sch_x=229 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14543 N$29085 N$29086 "Straight Waveguide" sch_x=229 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14544 N$29087 N$29088 "Straight Waveguide" sch_x=229 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14545 N$29089 N$29090 "Straight Waveguide" sch_x=229 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14546 N$29091 N$29092 "Straight Waveguide" sch_x=229 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14547 N$29093 N$29094 "Straight Waveguide" sch_x=229 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14548 N$29095 N$29096 "Straight Waveguide" sch_x=229 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14549 N$29097 N$29098 "Straight Waveguide" sch_x=229 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14550 N$29099 N$29100 "Straight Waveguide" sch_x=229 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14551 N$29101 N$29102 "Straight Waveguide" sch_x=229 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14552 N$29103 N$29104 "Straight Waveguide" sch_x=229 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14553 N$29105 N$29106 "Straight Waveguide" sch_x=229 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14554 N$29107 N$29108 "Straight Waveguide" sch_x=229 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14555 N$29109 N$29110 "Straight Waveguide" sch_x=229 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14556 N$29111 N$29112 "Straight Waveguide" sch_x=229 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14557 N$29113 N$29114 "Straight Waveguide" sch_x=229 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14558 N$29115 N$29116 "Straight Waveguide" sch_x=229 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14559 N$29117 N$29118 "Straight Waveguide" sch_x=229 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14560 N$29119 N$29120 "Straight Waveguide" sch_x=229 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14561 N$29121 N$29122 "Straight Waveguide" sch_x=229 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14562 N$29123 N$29124 "Straight Waveguide" sch_x=229 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14563 N$29125 N$29126 "Straight Waveguide" sch_x=229 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14564 N$29127 N$29128 "Straight Waveguide" sch_x=229 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14565 N$29129 N$29130 "Straight Waveguide" sch_x=229 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14566 N$29131 N$29132 "Straight Waveguide" sch_x=229 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14567 N$29133 N$29134 "Straight Waveguide" sch_x=229 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14568 N$29135 N$29136 "Straight Waveguide" sch_x=229 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14569 N$29137 N$29138 "Straight Waveguide" sch_x=229 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14570 N$29139 N$29140 "Straight Waveguide" sch_x=229 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14571 N$29141 N$29142 "Straight Waveguide" sch_x=229 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14572 N$29143 N$29144 "Straight Waveguide" sch_x=229 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14573 N$29145 N$29146 "Straight Waveguide" sch_x=229 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14574 N$29147 N$29148 "Straight Waveguide" sch_x=229 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14575 N$29149 N$29150 "Straight Waveguide" sch_x=229 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14576 N$29151 N$29152 "Straight Waveguide" sch_x=229 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14577 N$29153 N$29154 "Straight Waveguide" sch_x=229 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14578 N$29155 N$29156 "Straight Waveguide" sch_x=229 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14579 N$29157 N$29158 "Straight Waveguide" sch_x=229 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14580 N$29159 N$29160 "Straight Waveguide" sch_x=229 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14581 N$29161 N$29162 "Straight Waveguide" sch_x=229 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14582 N$29163 N$29164 "Straight Waveguide" sch_x=229 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14583 N$29165 N$29166 "Straight Waveguide" sch_x=229 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14584 N$29167 N$29168 "Straight Waveguide" sch_x=229 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14585 N$29169 N$29170 "Straight Waveguide" sch_x=229 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14586 N$29171 N$29172 "Straight Waveguide" sch_x=229 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14587 N$29173 N$29174 "Straight Waveguide" sch_x=229 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14588 N$29175 N$29176 "Straight Waveguide" sch_x=229 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14589 N$29177 N$29178 "Straight Waveguide" sch_x=229 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14590 N$29179 N$29180 "Straight Waveguide" sch_x=229 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14591 N$29181 N$29182 "Straight Waveguide" sch_x=229 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14592 N$29183 N$29184 "Straight Waveguide" sch_x=229 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14593 N$29185 N$29186 "Straight Waveguide" sch_x=229 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14594 N$29187 N$29188 "Straight Waveguide" sch_x=229 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14595 N$29189 N$29190 "Straight Waveguide" sch_x=229 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14596 N$29191 N$29192 "Straight Waveguide" sch_x=229 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14597 N$29193 N$29194 "Straight Waveguide" sch_x=229 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14598 N$29195 N$29196 "Straight Waveguide" sch_x=229 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14599 N$29197 N$29198 "Straight Waveguide" sch_x=229 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14600 N$29199 N$29200 "Straight Waveguide" sch_x=229 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14601 N$29201 N$29202 "Straight Waveguide" sch_x=229 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14602 N$29203 N$29204 "Straight Waveguide" sch_x=229 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14603 N$29205 N$29206 "Straight Waveguide" sch_x=227 sch_y=49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14604 N$29207 N$29208 "Straight Waveguide" sch_x=227 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14605 N$29209 N$29210 "Straight Waveguide" sch_x=227 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14606 N$29211 N$29212 "Straight Waveguide" sch_x=227 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14607 N$29213 N$29214 "Straight Waveguide" sch_x=227 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14608 N$29215 N$29216 "Straight Waveguide" sch_x=227 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14609 N$29217 N$29218 "Straight Waveguide" sch_x=227 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14610 N$29219 N$29220 "Straight Waveguide" sch_x=227 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14611 N$29221 N$29222 "Straight Waveguide" sch_x=227 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14612 N$29223 N$29224 "Straight Waveguide" sch_x=227 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14613 N$29225 N$29226 "Straight Waveguide" sch_x=227 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14614 N$29227 N$29228 "Straight Waveguide" sch_x=227 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14615 N$29229 N$29230 "Straight Waveguide" sch_x=227 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14616 N$29231 N$29232 "Straight Waveguide" sch_x=227 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14617 N$29233 N$29234 "Straight Waveguide" sch_x=227 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14618 N$29235 N$29236 "Straight Waveguide" sch_x=227 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14619 N$29237 N$29238 "Straight Waveguide" sch_x=227 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14620 N$29239 N$29240 "Straight Waveguide" sch_x=227 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14621 N$29241 N$29242 "Straight Waveguide" sch_x=227 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14622 N$29243 N$29244 "Straight Waveguide" sch_x=227 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14623 N$29245 N$29246 "Straight Waveguide" sch_x=227 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14624 N$29247 N$29248 "Straight Waveguide" sch_x=227 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14625 N$29249 N$29250 "Straight Waveguide" sch_x=227 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14626 N$29251 N$29252 "Straight Waveguide" sch_x=227 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14627 N$29253 N$29254 "Straight Waveguide" sch_x=227 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14628 N$29255 N$29256 "Straight Waveguide" sch_x=227 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14629 N$29257 N$29258 "Straight Waveguide" sch_x=227 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14630 N$29259 N$29260 "Straight Waveguide" sch_x=227 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14631 N$29261 N$29262 "Straight Waveguide" sch_x=227 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14632 N$29263 N$29264 "Straight Waveguide" sch_x=227 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14633 N$29265 N$29266 "Straight Waveguide" sch_x=227 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14634 N$29267 N$29268 "Straight Waveguide" sch_x=227 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14635 N$29269 N$29270 "Straight Waveguide" sch_x=227 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14636 N$29271 N$29272 "Straight Waveguide" sch_x=227 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14637 N$29273 N$29274 "Straight Waveguide" sch_x=227 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14638 N$29275 N$29276 "Straight Waveguide" sch_x=227 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14639 N$29277 N$29278 "Straight Waveguide" sch_x=227 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14640 N$29279 N$29280 "Straight Waveguide" sch_x=227 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14641 N$29281 N$29282 "Straight Waveguide" sch_x=227 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14642 N$29283 N$29284 "Straight Waveguide" sch_x=227 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14643 N$29285 N$29286 "Straight Waveguide" sch_x=227 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14644 N$29287 N$29288 "Straight Waveguide" sch_x=227 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14645 N$29289 N$29290 "Straight Waveguide" sch_x=227 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14646 N$29291 N$29292 "Straight Waveguide" sch_x=227 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14647 N$29293 N$29294 "Straight Waveguide" sch_x=227 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14648 N$29295 N$29296 "Straight Waveguide" sch_x=227 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14649 N$29297 N$29298 "Straight Waveguide" sch_x=227 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14650 N$29299 N$29300 "Straight Waveguide" sch_x=227 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14651 N$29301 N$29302 "Straight Waveguide" sch_x=227 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14652 N$29303 N$29304 "Straight Waveguide" sch_x=227 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14653 N$29305 N$29306 "Straight Waveguide" sch_x=227 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14654 N$29307 N$29308 "Straight Waveguide" sch_x=227 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14655 N$29309 N$29310 "Straight Waveguide" sch_x=227 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14656 N$29311 N$29312 "Straight Waveguide" sch_x=227 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14657 N$29313 N$29314 "Straight Waveguide" sch_x=227 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14658 N$29315 N$29316 "Straight Waveguide" sch_x=227 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14659 N$29317 N$29318 "Straight Waveguide" sch_x=227 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14660 N$29319 N$29320 "Straight Waveguide" sch_x=227 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14661 N$29321 N$29322 "Straight Waveguide" sch_x=227 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14662 N$29323 N$29324 "Straight Waveguide" sch_x=227 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14663 N$29325 N$29326 "Straight Waveguide" sch_x=227 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14664 N$29327 N$29328 "Straight Waveguide" sch_x=227 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14665 N$29329 N$29330 "Straight Waveguide" sch_x=227 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14666 N$29331 N$29332 "Straight Waveguide" sch_x=227 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14667 N$29333 N$29334 "Straight Waveguide" sch_x=227 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14668 N$29335 N$29336 "Straight Waveguide" sch_x=227 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14669 N$29337 N$29338 "Straight Waveguide" sch_x=227 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14670 N$29339 N$29340 "Straight Waveguide" sch_x=227 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14671 N$29341 N$29342 "Straight Waveguide" sch_x=227 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14672 N$29343 N$29344 "Straight Waveguide" sch_x=227 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14673 N$29345 N$29346 "Straight Waveguide" sch_x=227 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14674 N$29347 N$29348 "Straight Waveguide" sch_x=227 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14675 N$29349 N$29350 "Straight Waveguide" sch_x=227 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14676 N$29351 N$29352 "Straight Waveguide" sch_x=227 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14677 N$29353 N$29354 "Straight Waveguide" sch_x=227 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14678 N$29355 N$29356 "Straight Waveguide" sch_x=227 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14679 N$29357 N$29358 "Straight Waveguide" sch_x=227 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14680 N$29359 N$29360 "Straight Waveguide" sch_x=227 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14681 N$29361 N$29362 "Straight Waveguide" sch_x=227 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14682 N$29363 N$29364 "Straight Waveguide" sch_x=227 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14683 N$29365 N$29366 "Straight Waveguide" sch_x=227 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14684 N$29367 N$29368 "Straight Waveguide" sch_x=227 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14685 N$29369 N$29370 "Straight Waveguide" sch_x=227 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14686 N$29371 N$29372 "Straight Waveguide" sch_x=227 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14687 N$29373 N$29374 "Straight Waveguide" sch_x=227 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14688 N$29375 N$29376 "Straight Waveguide" sch_x=227 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14689 N$29377 N$29378 "Straight Waveguide" sch_x=227 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14690 N$29379 N$29380 "Straight Waveguide" sch_x=227 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14691 N$29381 N$29382 "Straight Waveguide" sch_x=227 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14692 N$29383 N$29384 "Straight Waveguide" sch_x=227 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14693 N$29385 N$29386 "Straight Waveguide" sch_x=227 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14694 N$29387 N$29388 "Straight Waveguide" sch_x=227 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14695 N$29389 N$29390 "Straight Waveguide" sch_x=227 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14696 N$29391 N$29392 "Straight Waveguide" sch_x=227 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14697 N$29393 N$29394 "Straight Waveguide" sch_x=227 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14698 N$29395 N$29396 "Straight Waveguide" sch_x=227 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14699 N$29397 N$29398 "Straight Waveguide" sch_x=227 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14700 N$29399 N$29400 "Straight Waveguide" sch_x=227 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14701 N$29401 N$29402 "Straight Waveguide" sch_x=227 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14702 N$29403 N$29404 "Straight Waveguide" sch_x=227 sch_y=-49.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14703 N$29405 N$29406 "Straight Waveguide" sch_x=225 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14704 N$29407 N$29408 "Straight Waveguide" sch_x=225 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14705 N$29409 N$29410 "Straight Waveguide" sch_x=225 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14706 N$29411 N$29412 "Straight Waveguide" sch_x=225 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14707 N$29413 N$29414 "Straight Waveguide" sch_x=225 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14708 N$29415 N$29416 "Straight Waveguide" sch_x=225 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14709 N$29417 N$29418 "Straight Waveguide" sch_x=225 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14710 N$29419 N$29420 "Straight Waveguide" sch_x=225 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14711 N$29421 N$29422 "Straight Waveguide" sch_x=225 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14712 N$29423 N$29424 "Straight Waveguide" sch_x=225 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14713 N$29425 N$29426 "Straight Waveguide" sch_x=225 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14714 N$29427 N$29428 "Straight Waveguide" sch_x=225 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14715 N$29429 N$29430 "Straight Waveguide" sch_x=225 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14716 N$29431 N$29432 "Straight Waveguide" sch_x=225 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14717 N$29433 N$29434 "Straight Waveguide" sch_x=225 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14718 N$29435 N$29436 "Straight Waveguide" sch_x=225 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14719 N$29437 N$29438 "Straight Waveguide" sch_x=225 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14720 N$29439 N$29440 "Straight Waveguide" sch_x=225 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14721 N$29441 N$29442 "Straight Waveguide" sch_x=225 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14722 N$29443 N$29444 "Straight Waveguide" sch_x=225 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14723 N$29445 N$29446 "Straight Waveguide" sch_x=225 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14724 N$29447 N$29448 "Straight Waveguide" sch_x=225 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14725 N$29449 N$29450 "Straight Waveguide" sch_x=225 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14726 N$29451 N$29452 "Straight Waveguide" sch_x=225 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14727 N$29453 N$29454 "Straight Waveguide" sch_x=225 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14728 N$29455 N$29456 "Straight Waveguide" sch_x=225 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14729 N$29457 N$29458 "Straight Waveguide" sch_x=225 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14730 N$29459 N$29460 "Straight Waveguide" sch_x=225 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14731 N$29461 N$29462 "Straight Waveguide" sch_x=225 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14732 N$29463 N$29464 "Straight Waveguide" sch_x=225 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14733 N$29465 N$29466 "Straight Waveguide" sch_x=225 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14734 N$29467 N$29468 "Straight Waveguide" sch_x=225 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14735 N$29469 N$29470 "Straight Waveguide" sch_x=225 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14736 N$29471 N$29472 "Straight Waveguide" sch_x=225 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14737 N$29473 N$29474 "Straight Waveguide" sch_x=225 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14738 N$29475 N$29476 "Straight Waveguide" sch_x=225 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14739 N$29477 N$29478 "Straight Waveguide" sch_x=225 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14740 N$29479 N$29480 "Straight Waveguide" sch_x=225 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14741 N$29481 N$29482 "Straight Waveguide" sch_x=225 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14742 N$29483 N$29484 "Straight Waveguide" sch_x=225 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14743 N$29485 N$29486 "Straight Waveguide" sch_x=225 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14744 N$29487 N$29488 "Straight Waveguide" sch_x=225 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14745 N$29489 N$29490 "Straight Waveguide" sch_x=225 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14746 N$29491 N$29492 "Straight Waveguide" sch_x=225 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14747 N$29493 N$29494 "Straight Waveguide" sch_x=225 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14748 N$29495 N$29496 "Straight Waveguide" sch_x=225 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14749 N$29497 N$29498 "Straight Waveguide" sch_x=225 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14750 N$29499 N$29500 "Straight Waveguide" sch_x=225 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14751 N$29501 N$29502 "Straight Waveguide" sch_x=225 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14752 N$29503 N$29504 "Straight Waveguide" sch_x=225 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14753 N$29505 N$29506 "Straight Waveguide" sch_x=225 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14754 N$29507 N$29508 "Straight Waveguide" sch_x=225 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14755 N$29509 N$29510 "Straight Waveguide" sch_x=225 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14756 N$29511 N$29512 "Straight Waveguide" sch_x=225 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14757 N$29513 N$29514 "Straight Waveguide" sch_x=225 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14758 N$29515 N$29516 "Straight Waveguide" sch_x=225 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14759 N$29517 N$29518 "Straight Waveguide" sch_x=225 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14760 N$29519 N$29520 "Straight Waveguide" sch_x=225 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14761 N$29521 N$29522 "Straight Waveguide" sch_x=225 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14762 N$29523 N$29524 "Straight Waveguide" sch_x=225 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14763 N$29525 N$29526 "Straight Waveguide" sch_x=225 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14764 N$29527 N$29528 "Straight Waveguide" sch_x=225 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14765 N$29529 N$29530 "Straight Waveguide" sch_x=225 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14766 N$29531 N$29532 "Straight Waveguide" sch_x=225 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14767 N$29533 N$29534 "Straight Waveguide" sch_x=225 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14768 N$29535 N$29536 "Straight Waveguide" sch_x=225 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14769 N$29537 N$29538 "Straight Waveguide" sch_x=225 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14770 N$29539 N$29540 "Straight Waveguide" sch_x=225 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14771 N$29541 N$29542 "Straight Waveguide" sch_x=225 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14772 N$29543 N$29544 "Straight Waveguide" sch_x=225 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14773 N$29545 N$29546 "Straight Waveguide" sch_x=225 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14774 N$29547 N$29548 "Straight Waveguide" sch_x=225 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14775 N$29549 N$29550 "Straight Waveguide" sch_x=225 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14776 N$29551 N$29552 "Straight Waveguide" sch_x=225 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14777 N$29553 N$29554 "Straight Waveguide" sch_x=225 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14778 N$29555 N$29556 "Straight Waveguide" sch_x=225 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14779 N$29557 N$29558 "Straight Waveguide" sch_x=225 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14780 N$29559 N$29560 "Straight Waveguide" sch_x=225 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14781 N$29561 N$29562 "Straight Waveguide" sch_x=225 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14782 N$29563 N$29564 "Straight Waveguide" sch_x=225 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14783 N$29565 N$29566 "Straight Waveguide" sch_x=225 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14784 N$29567 N$29568 "Straight Waveguide" sch_x=225 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14785 N$29569 N$29570 "Straight Waveguide" sch_x=225 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14786 N$29571 N$29572 "Straight Waveguide" sch_x=225 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14787 N$29573 N$29574 "Straight Waveguide" sch_x=225 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14788 N$29575 N$29576 "Straight Waveguide" sch_x=225 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14789 N$29577 N$29578 "Straight Waveguide" sch_x=225 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14790 N$29579 N$29580 "Straight Waveguide" sch_x=225 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14791 N$29581 N$29582 "Straight Waveguide" sch_x=225 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14792 N$29583 N$29584 "Straight Waveguide" sch_x=225 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14793 N$29585 N$29586 "Straight Waveguide" sch_x=225 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14794 N$29587 N$29588 "Straight Waveguide" sch_x=225 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14795 N$29589 N$29590 "Straight Waveguide" sch_x=225 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14796 N$29591 N$29592 "Straight Waveguide" sch_x=225 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14797 N$29593 N$29594 "Straight Waveguide" sch_x=225 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14798 N$29595 N$29596 "Straight Waveguide" sch_x=225 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14799 N$29597 N$29598 "Straight Waveguide" sch_x=225 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14800 N$29599 N$29600 "Straight Waveguide" sch_x=225 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14801 N$29601 N$29602 "Straight Waveguide" sch_x=223 sch_y=47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14802 N$29603 N$29604 "Straight Waveguide" sch_x=223 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14803 N$29605 N$29606 "Straight Waveguide" sch_x=223 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14804 N$29607 N$29608 "Straight Waveguide" sch_x=223 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14805 N$29609 N$29610 "Straight Waveguide" sch_x=223 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14806 N$29611 N$29612 "Straight Waveguide" sch_x=223 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14807 N$29613 N$29614 "Straight Waveguide" sch_x=223 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14808 N$29615 N$29616 "Straight Waveguide" sch_x=223 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14809 N$29617 N$29618 "Straight Waveguide" sch_x=223 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14810 N$29619 N$29620 "Straight Waveguide" sch_x=223 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14811 N$29621 N$29622 "Straight Waveguide" sch_x=223 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14812 N$29623 N$29624 "Straight Waveguide" sch_x=223 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14813 N$29625 N$29626 "Straight Waveguide" sch_x=223 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14814 N$29627 N$29628 "Straight Waveguide" sch_x=223 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14815 N$29629 N$29630 "Straight Waveguide" sch_x=223 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14816 N$29631 N$29632 "Straight Waveguide" sch_x=223 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14817 N$29633 N$29634 "Straight Waveguide" sch_x=223 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14818 N$29635 N$29636 "Straight Waveguide" sch_x=223 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14819 N$29637 N$29638 "Straight Waveguide" sch_x=223 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14820 N$29639 N$29640 "Straight Waveguide" sch_x=223 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14821 N$29641 N$29642 "Straight Waveguide" sch_x=223 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14822 N$29643 N$29644 "Straight Waveguide" sch_x=223 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14823 N$29645 N$29646 "Straight Waveguide" sch_x=223 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14824 N$29647 N$29648 "Straight Waveguide" sch_x=223 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14825 N$29649 N$29650 "Straight Waveguide" sch_x=223 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14826 N$29651 N$29652 "Straight Waveguide" sch_x=223 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14827 N$29653 N$29654 "Straight Waveguide" sch_x=223 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14828 N$29655 N$29656 "Straight Waveguide" sch_x=223 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14829 N$29657 N$29658 "Straight Waveguide" sch_x=223 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14830 N$29659 N$29660 "Straight Waveguide" sch_x=223 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14831 N$29661 N$29662 "Straight Waveguide" sch_x=223 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14832 N$29663 N$29664 "Straight Waveguide" sch_x=223 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14833 N$29665 N$29666 "Straight Waveguide" sch_x=223 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14834 N$29667 N$29668 "Straight Waveguide" sch_x=223 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14835 N$29669 N$29670 "Straight Waveguide" sch_x=223 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14836 N$29671 N$29672 "Straight Waveguide" sch_x=223 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14837 N$29673 N$29674 "Straight Waveguide" sch_x=223 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14838 N$29675 N$29676 "Straight Waveguide" sch_x=223 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14839 N$29677 N$29678 "Straight Waveguide" sch_x=223 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14840 N$29679 N$29680 "Straight Waveguide" sch_x=223 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14841 N$29681 N$29682 "Straight Waveguide" sch_x=223 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14842 N$29683 N$29684 "Straight Waveguide" sch_x=223 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14843 N$29685 N$29686 "Straight Waveguide" sch_x=223 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14844 N$29687 N$29688 "Straight Waveguide" sch_x=223 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14845 N$29689 N$29690 "Straight Waveguide" sch_x=223 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14846 N$29691 N$29692 "Straight Waveguide" sch_x=223 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14847 N$29693 N$29694 "Straight Waveguide" sch_x=223 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14848 N$29695 N$29696 "Straight Waveguide" sch_x=223 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14849 N$29697 N$29698 "Straight Waveguide" sch_x=223 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14850 N$29699 N$29700 "Straight Waveguide" sch_x=223 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14851 N$29701 N$29702 "Straight Waveguide" sch_x=223 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14852 N$29703 N$29704 "Straight Waveguide" sch_x=223 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14853 N$29705 N$29706 "Straight Waveguide" sch_x=223 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14854 N$29707 N$29708 "Straight Waveguide" sch_x=223 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14855 N$29709 N$29710 "Straight Waveguide" sch_x=223 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14856 N$29711 N$29712 "Straight Waveguide" sch_x=223 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14857 N$29713 N$29714 "Straight Waveguide" sch_x=223 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14858 N$29715 N$29716 "Straight Waveguide" sch_x=223 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14859 N$29717 N$29718 "Straight Waveguide" sch_x=223 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14860 N$29719 N$29720 "Straight Waveguide" sch_x=223 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14861 N$29721 N$29722 "Straight Waveguide" sch_x=223 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14862 N$29723 N$29724 "Straight Waveguide" sch_x=223 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14863 N$29725 N$29726 "Straight Waveguide" sch_x=223 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14864 N$29727 N$29728 "Straight Waveguide" sch_x=223 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14865 N$29729 N$29730 "Straight Waveguide" sch_x=223 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14866 N$29731 N$29732 "Straight Waveguide" sch_x=223 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14867 N$29733 N$29734 "Straight Waveguide" sch_x=223 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14868 N$29735 N$29736 "Straight Waveguide" sch_x=223 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14869 N$29737 N$29738 "Straight Waveguide" sch_x=223 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14870 N$29739 N$29740 "Straight Waveguide" sch_x=223 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14871 N$29741 N$29742 "Straight Waveguide" sch_x=223 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14872 N$29743 N$29744 "Straight Waveguide" sch_x=223 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14873 N$29745 N$29746 "Straight Waveguide" sch_x=223 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14874 N$29747 N$29748 "Straight Waveguide" sch_x=223 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14875 N$29749 N$29750 "Straight Waveguide" sch_x=223 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14876 N$29751 N$29752 "Straight Waveguide" sch_x=223 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14877 N$29753 N$29754 "Straight Waveguide" sch_x=223 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14878 N$29755 N$29756 "Straight Waveguide" sch_x=223 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14879 N$29757 N$29758 "Straight Waveguide" sch_x=223 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14880 N$29759 N$29760 "Straight Waveguide" sch_x=223 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14881 N$29761 N$29762 "Straight Waveguide" sch_x=223 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14882 N$29763 N$29764 "Straight Waveguide" sch_x=223 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14883 N$29765 N$29766 "Straight Waveguide" sch_x=223 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14884 N$29767 N$29768 "Straight Waveguide" sch_x=223 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14885 N$29769 N$29770 "Straight Waveguide" sch_x=223 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14886 N$29771 N$29772 "Straight Waveguide" sch_x=223 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14887 N$29773 N$29774 "Straight Waveguide" sch_x=223 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14888 N$29775 N$29776 "Straight Waveguide" sch_x=223 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14889 N$29777 N$29778 "Straight Waveguide" sch_x=223 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14890 N$29779 N$29780 "Straight Waveguide" sch_x=223 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14891 N$29781 N$29782 "Straight Waveguide" sch_x=223 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14892 N$29783 N$29784 "Straight Waveguide" sch_x=223 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14893 N$29785 N$29786 "Straight Waveguide" sch_x=223 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14894 N$29787 N$29788 "Straight Waveguide" sch_x=223 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14895 N$29789 N$29790 "Straight Waveguide" sch_x=223 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14896 N$29791 N$29792 "Straight Waveguide" sch_x=223 sch_y=-47.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14897 N$29793 N$29794 "Straight Waveguide" sch_x=221 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14898 N$29795 N$29796 "Straight Waveguide" sch_x=221 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14899 N$29797 N$29798 "Straight Waveguide" sch_x=221 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14900 N$29799 N$29800 "Straight Waveguide" sch_x=221 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14901 N$29801 N$29802 "Straight Waveguide" sch_x=221 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14902 N$29803 N$29804 "Straight Waveguide" sch_x=221 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14903 N$29805 N$29806 "Straight Waveguide" sch_x=221 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14904 N$29807 N$29808 "Straight Waveguide" sch_x=221 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14905 N$29809 N$29810 "Straight Waveguide" sch_x=221 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14906 N$29811 N$29812 "Straight Waveguide" sch_x=221 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14907 N$29813 N$29814 "Straight Waveguide" sch_x=221 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14908 N$29815 N$29816 "Straight Waveguide" sch_x=221 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14909 N$29817 N$29818 "Straight Waveguide" sch_x=221 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14910 N$29819 N$29820 "Straight Waveguide" sch_x=221 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14911 N$29821 N$29822 "Straight Waveguide" sch_x=221 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14912 N$29823 N$29824 "Straight Waveguide" sch_x=221 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14913 N$29825 N$29826 "Straight Waveguide" sch_x=221 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14914 N$29827 N$29828 "Straight Waveguide" sch_x=221 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14915 N$29829 N$29830 "Straight Waveguide" sch_x=221 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14916 N$29831 N$29832 "Straight Waveguide" sch_x=221 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14917 N$29833 N$29834 "Straight Waveguide" sch_x=221 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14918 N$29835 N$29836 "Straight Waveguide" sch_x=221 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14919 N$29837 N$29838 "Straight Waveguide" sch_x=221 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14920 N$29839 N$29840 "Straight Waveguide" sch_x=221 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14921 N$29841 N$29842 "Straight Waveguide" sch_x=221 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14922 N$29843 N$29844 "Straight Waveguide" sch_x=221 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14923 N$29845 N$29846 "Straight Waveguide" sch_x=221 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14924 N$29847 N$29848 "Straight Waveguide" sch_x=221 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14925 N$29849 N$29850 "Straight Waveguide" sch_x=221 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14926 N$29851 N$29852 "Straight Waveguide" sch_x=221 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14927 N$29853 N$29854 "Straight Waveguide" sch_x=221 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14928 N$29855 N$29856 "Straight Waveguide" sch_x=221 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14929 N$29857 N$29858 "Straight Waveguide" sch_x=221 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14930 N$29859 N$29860 "Straight Waveguide" sch_x=221 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14931 N$29861 N$29862 "Straight Waveguide" sch_x=221 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14932 N$29863 N$29864 "Straight Waveguide" sch_x=221 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14933 N$29865 N$29866 "Straight Waveguide" sch_x=221 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14934 N$29867 N$29868 "Straight Waveguide" sch_x=221 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14935 N$29869 N$29870 "Straight Waveguide" sch_x=221 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14936 N$29871 N$29872 "Straight Waveguide" sch_x=221 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14937 N$29873 N$29874 "Straight Waveguide" sch_x=221 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14938 N$29875 N$29876 "Straight Waveguide" sch_x=221 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14939 N$29877 N$29878 "Straight Waveguide" sch_x=221 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14940 N$29879 N$29880 "Straight Waveguide" sch_x=221 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14941 N$29881 N$29882 "Straight Waveguide" sch_x=221 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14942 N$29883 N$29884 "Straight Waveguide" sch_x=221 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14943 N$29885 N$29886 "Straight Waveguide" sch_x=221 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14944 N$29887 N$29888 "Straight Waveguide" sch_x=221 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14945 N$29889 N$29890 "Straight Waveguide" sch_x=221 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14946 N$29891 N$29892 "Straight Waveguide" sch_x=221 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14947 N$29893 N$29894 "Straight Waveguide" sch_x=221 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14948 N$29895 N$29896 "Straight Waveguide" sch_x=221 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14949 N$29897 N$29898 "Straight Waveguide" sch_x=221 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14950 N$29899 N$29900 "Straight Waveguide" sch_x=221 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14951 N$29901 N$29902 "Straight Waveguide" sch_x=221 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14952 N$29903 N$29904 "Straight Waveguide" sch_x=221 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14953 N$29905 N$29906 "Straight Waveguide" sch_x=221 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14954 N$29907 N$29908 "Straight Waveguide" sch_x=221 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14955 N$29909 N$29910 "Straight Waveguide" sch_x=221 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14956 N$29911 N$29912 "Straight Waveguide" sch_x=221 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14957 N$29913 N$29914 "Straight Waveguide" sch_x=221 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14958 N$29915 N$29916 "Straight Waveguide" sch_x=221 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14959 N$29917 N$29918 "Straight Waveguide" sch_x=221 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14960 N$29919 N$29920 "Straight Waveguide" sch_x=221 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14961 N$29921 N$29922 "Straight Waveguide" sch_x=221 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14962 N$29923 N$29924 "Straight Waveguide" sch_x=221 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14963 N$29925 N$29926 "Straight Waveguide" sch_x=221 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14964 N$29927 N$29928 "Straight Waveguide" sch_x=221 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14965 N$29929 N$29930 "Straight Waveguide" sch_x=221 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14966 N$29931 N$29932 "Straight Waveguide" sch_x=221 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14967 N$29933 N$29934 "Straight Waveguide" sch_x=221 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14968 N$29935 N$29936 "Straight Waveguide" sch_x=221 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14969 N$29937 N$29938 "Straight Waveguide" sch_x=221 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14970 N$29939 N$29940 "Straight Waveguide" sch_x=221 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14971 N$29941 N$29942 "Straight Waveguide" sch_x=221 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14972 N$29943 N$29944 "Straight Waveguide" sch_x=221 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14973 N$29945 N$29946 "Straight Waveguide" sch_x=221 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14974 N$29947 N$29948 "Straight Waveguide" sch_x=221 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14975 N$29949 N$29950 "Straight Waveguide" sch_x=221 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14976 N$29951 N$29952 "Straight Waveguide" sch_x=221 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14977 N$29953 N$29954 "Straight Waveguide" sch_x=221 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14978 N$29955 N$29956 "Straight Waveguide" sch_x=221 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14979 N$29957 N$29958 "Straight Waveguide" sch_x=221 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14980 N$29959 N$29960 "Straight Waveguide" sch_x=221 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14981 N$29961 N$29962 "Straight Waveguide" sch_x=221 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14982 N$29963 N$29964 "Straight Waveguide" sch_x=221 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14983 N$29965 N$29966 "Straight Waveguide" sch_x=221 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14984 N$29967 N$29968 "Straight Waveguide" sch_x=221 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14985 N$29969 N$29970 "Straight Waveguide" sch_x=221 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14986 N$29971 N$29972 "Straight Waveguide" sch_x=221 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14987 N$29973 N$29974 "Straight Waveguide" sch_x=221 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14988 N$29975 N$29976 "Straight Waveguide" sch_x=221 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14989 N$29977 N$29978 "Straight Waveguide" sch_x=221 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14990 N$29979 N$29980 "Straight Waveguide" sch_x=221 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14991 N$29981 N$29982 "Straight Waveguide" sch_x=219 sch_y=45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14992 N$29983 N$29984 "Straight Waveguide" sch_x=219 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14993 N$29985 N$29986 "Straight Waveguide" sch_x=219 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14994 N$29987 N$29988 "Straight Waveguide" sch_x=219 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14995 N$29989 N$29990 "Straight Waveguide" sch_x=219 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14996 N$29991 N$29992 "Straight Waveguide" sch_x=219 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14997 N$29993 N$29994 "Straight Waveguide" sch_x=219 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14998 N$29995 N$29996 "Straight Waveguide" sch_x=219 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14999 N$29997 N$29998 "Straight Waveguide" sch_x=219 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15000 N$29999 N$30000 "Straight Waveguide" sch_x=219 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15001 N$30001 N$30002 "Straight Waveguide" sch_x=219 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15002 N$30003 N$30004 "Straight Waveguide" sch_x=219 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15003 N$30005 N$30006 "Straight Waveguide" sch_x=219 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15004 N$30007 N$30008 "Straight Waveguide" sch_x=219 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15005 N$30009 N$30010 "Straight Waveguide" sch_x=219 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15006 N$30011 N$30012 "Straight Waveguide" sch_x=219 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15007 N$30013 N$30014 "Straight Waveguide" sch_x=219 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15008 N$30015 N$30016 "Straight Waveguide" sch_x=219 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15009 N$30017 N$30018 "Straight Waveguide" sch_x=219 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15010 N$30019 N$30020 "Straight Waveguide" sch_x=219 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15011 N$30021 N$30022 "Straight Waveguide" sch_x=219 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15012 N$30023 N$30024 "Straight Waveguide" sch_x=219 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15013 N$30025 N$30026 "Straight Waveguide" sch_x=219 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15014 N$30027 N$30028 "Straight Waveguide" sch_x=219 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15015 N$30029 N$30030 "Straight Waveguide" sch_x=219 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15016 N$30031 N$30032 "Straight Waveguide" sch_x=219 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15017 N$30033 N$30034 "Straight Waveguide" sch_x=219 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15018 N$30035 N$30036 "Straight Waveguide" sch_x=219 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15019 N$30037 N$30038 "Straight Waveguide" sch_x=219 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15020 N$30039 N$30040 "Straight Waveguide" sch_x=219 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15021 N$30041 N$30042 "Straight Waveguide" sch_x=219 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15022 N$30043 N$30044 "Straight Waveguide" sch_x=219 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15023 N$30045 N$30046 "Straight Waveguide" sch_x=219 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15024 N$30047 N$30048 "Straight Waveguide" sch_x=219 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15025 N$30049 N$30050 "Straight Waveguide" sch_x=219 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15026 N$30051 N$30052 "Straight Waveguide" sch_x=219 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15027 N$30053 N$30054 "Straight Waveguide" sch_x=219 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15028 N$30055 N$30056 "Straight Waveguide" sch_x=219 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15029 N$30057 N$30058 "Straight Waveguide" sch_x=219 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15030 N$30059 N$30060 "Straight Waveguide" sch_x=219 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15031 N$30061 N$30062 "Straight Waveguide" sch_x=219 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15032 N$30063 N$30064 "Straight Waveguide" sch_x=219 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15033 N$30065 N$30066 "Straight Waveguide" sch_x=219 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15034 N$30067 N$30068 "Straight Waveguide" sch_x=219 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15035 N$30069 N$30070 "Straight Waveguide" sch_x=219 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15036 N$30071 N$30072 "Straight Waveguide" sch_x=219 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15037 N$30073 N$30074 "Straight Waveguide" sch_x=219 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15038 N$30075 N$30076 "Straight Waveguide" sch_x=219 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15039 N$30077 N$30078 "Straight Waveguide" sch_x=219 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15040 N$30079 N$30080 "Straight Waveguide" sch_x=219 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15041 N$30081 N$30082 "Straight Waveguide" sch_x=219 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15042 N$30083 N$30084 "Straight Waveguide" sch_x=219 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15043 N$30085 N$30086 "Straight Waveguide" sch_x=219 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15044 N$30087 N$30088 "Straight Waveguide" sch_x=219 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15045 N$30089 N$30090 "Straight Waveguide" sch_x=219 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15046 N$30091 N$30092 "Straight Waveguide" sch_x=219 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15047 N$30093 N$30094 "Straight Waveguide" sch_x=219 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15048 N$30095 N$30096 "Straight Waveguide" sch_x=219 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15049 N$30097 N$30098 "Straight Waveguide" sch_x=219 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15050 N$30099 N$30100 "Straight Waveguide" sch_x=219 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15051 N$30101 N$30102 "Straight Waveguide" sch_x=219 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15052 N$30103 N$30104 "Straight Waveguide" sch_x=219 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15053 N$30105 N$30106 "Straight Waveguide" sch_x=219 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15054 N$30107 N$30108 "Straight Waveguide" sch_x=219 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15055 N$30109 N$30110 "Straight Waveguide" sch_x=219 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15056 N$30111 N$30112 "Straight Waveguide" sch_x=219 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15057 N$30113 N$30114 "Straight Waveguide" sch_x=219 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15058 N$30115 N$30116 "Straight Waveguide" sch_x=219 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15059 N$30117 N$30118 "Straight Waveguide" sch_x=219 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15060 N$30119 N$30120 "Straight Waveguide" sch_x=219 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15061 N$30121 N$30122 "Straight Waveguide" sch_x=219 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15062 N$30123 N$30124 "Straight Waveguide" sch_x=219 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15063 N$30125 N$30126 "Straight Waveguide" sch_x=219 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15064 N$30127 N$30128 "Straight Waveguide" sch_x=219 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15065 N$30129 N$30130 "Straight Waveguide" sch_x=219 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15066 N$30131 N$30132 "Straight Waveguide" sch_x=219 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15067 N$30133 N$30134 "Straight Waveguide" sch_x=219 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15068 N$30135 N$30136 "Straight Waveguide" sch_x=219 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15069 N$30137 N$30138 "Straight Waveguide" sch_x=219 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15070 N$30139 N$30140 "Straight Waveguide" sch_x=219 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15071 N$30141 N$30142 "Straight Waveguide" sch_x=219 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15072 N$30143 N$30144 "Straight Waveguide" sch_x=219 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15073 N$30145 N$30146 "Straight Waveguide" sch_x=219 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15074 N$30147 N$30148 "Straight Waveguide" sch_x=219 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15075 N$30149 N$30150 "Straight Waveguide" sch_x=219 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15076 N$30151 N$30152 "Straight Waveguide" sch_x=219 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15077 N$30153 N$30154 "Straight Waveguide" sch_x=219 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15078 N$30155 N$30156 "Straight Waveguide" sch_x=219 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15079 N$30157 N$30158 "Straight Waveguide" sch_x=219 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15080 N$30159 N$30160 "Straight Waveguide" sch_x=219 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15081 N$30161 N$30162 "Straight Waveguide" sch_x=219 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15082 N$30163 N$30164 "Straight Waveguide" sch_x=219 sch_y=-45.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15083 N$30165 N$30166 "Straight Waveguide" sch_x=217 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15084 N$30167 N$30168 "Straight Waveguide" sch_x=217 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15085 N$30169 N$30170 "Straight Waveguide" sch_x=217 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15086 N$30171 N$30172 "Straight Waveguide" sch_x=217 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15087 N$30173 N$30174 "Straight Waveguide" sch_x=217 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15088 N$30175 N$30176 "Straight Waveguide" sch_x=217 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15089 N$30177 N$30178 "Straight Waveguide" sch_x=217 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15090 N$30179 N$30180 "Straight Waveguide" sch_x=217 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15091 N$30181 N$30182 "Straight Waveguide" sch_x=217 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15092 N$30183 N$30184 "Straight Waveguide" sch_x=217 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15093 N$30185 N$30186 "Straight Waveguide" sch_x=217 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15094 N$30187 N$30188 "Straight Waveguide" sch_x=217 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15095 N$30189 N$30190 "Straight Waveguide" sch_x=217 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15096 N$30191 N$30192 "Straight Waveguide" sch_x=217 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15097 N$30193 N$30194 "Straight Waveguide" sch_x=217 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15098 N$30195 N$30196 "Straight Waveguide" sch_x=217 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15099 N$30197 N$30198 "Straight Waveguide" sch_x=217 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15100 N$30199 N$30200 "Straight Waveguide" sch_x=217 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15101 N$30201 N$30202 "Straight Waveguide" sch_x=217 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15102 N$30203 N$30204 "Straight Waveguide" sch_x=217 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15103 N$30205 N$30206 "Straight Waveguide" sch_x=217 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15104 N$30207 N$30208 "Straight Waveguide" sch_x=217 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15105 N$30209 N$30210 "Straight Waveguide" sch_x=217 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15106 N$30211 N$30212 "Straight Waveguide" sch_x=217 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15107 N$30213 N$30214 "Straight Waveguide" sch_x=217 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15108 N$30215 N$30216 "Straight Waveguide" sch_x=217 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15109 N$30217 N$30218 "Straight Waveguide" sch_x=217 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15110 N$30219 N$30220 "Straight Waveguide" sch_x=217 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15111 N$30221 N$30222 "Straight Waveguide" sch_x=217 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15112 N$30223 N$30224 "Straight Waveguide" sch_x=217 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15113 N$30225 N$30226 "Straight Waveguide" sch_x=217 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15114 N$30227 N$30228 "Straight Waveguide" sch_x=217 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15115 N$30229 N$30230 "Straight Waveguide" sch_x=217 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15116 N$30231 N$30232 "Straight Waveguide" sch_x=217 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15117 N$30233 N$30234 "Straight Waveguide" sch_x=217 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15118 N$30235 N$30236 "Straight Waveguide" sch_x=217 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15119 N$30237 N$30238 "Straight Waveguide" sch_x=217 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15120 N$30239 N$30240 "Straight Waveguide" sch_x=217 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15121 N$30241 N$30242 "Straight Waveguide" sch_x=217 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15122 N$30243 N$30244 "Straight Waveguide" sch_x=217 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15123 N$30245 N$30246 "Straight Waveguide" sch_x=217 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15124 N$30247 N$30248 "Straight Waveguide" sch_x=217 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15125 N$30249 N$30250 "Straight Waveguide" sch_x=217 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15126 N$30251 N$30252 "Straight Waveguide" sch_x=217 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15127 N$30253 N$30254 "Straight Waveguide" sch_x=217 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15128 N$30255 N$30256 "Straight Waveguide" sch_x=217 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15129 N$30257 N$30258 "Straight Waveguide" sch_x=217 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15130 N$30259 N$30260 "Straight Waveguide" sch_x=217 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15131 N$30261 N$30262 "Straight Waveguide" sch_x=217 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15132 N$30263 N$30264 "Straight Waveguide" sch_x=217 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15133 N$30265 N$30266 "Straight Waveguide" sch_x=217 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15134 N$30267 N$30268 "Straight Waveguide" sch_x=217 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15135 N$30269 N$30270 "Straight Waveguide" sch_x=217 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15136 N$30271 N$30272 "Straight Waveguide" sch_x=217 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15137 N$30273 N$30274 "Straight Waveguide" sch_x=217 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15138 N$30275 N$30276 "Straight Waveguide" sch_x=217 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15139 N$30277 N$30278 "Straight Waveguide" sch_x=217 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15140 N$30279 N$30280 "Straight Waveguide" sch_x=217 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15141 N$30281 N$30282 "Straight Waveguide" sch_x=217 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15142 N$30283 N$30284 "Straight Waveguide" sch_x=217 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15143 N$30285 N$30286 "Straight Waveguide" sch_x=217 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15144 N$30287 N$30288 "Straight Waveguide" sch_x=217 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15145 N$30289 N$30290 "Straight Waveguide" sch_x=217 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15146 N$30291 N$30292 "Straight Waveguide" sch_x=217 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15147 N$30293 N$30294 "Straight Waveguide" sch_x=217 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15148 N$30295 N$30296 "Straight Waveguide" sch_x=217 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15149 N$30297 N$30298 "Straight Waveguide" sch_x=217 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15150 N$30299 N$30300 "Straight Waveguide" sch_x=217 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15151 N$30301 N$30302 "Straight Waveguide" sch_x=217 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15152 N$30303 N$30304 "Straight Waveguide" sch_x=217 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15153 N$30305 N$30306 "Straight Waveguide" sch_x=217 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15154 N$30307 N$30308 "Straight Waveguide" sch_x=217 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15155 N$30309 N$30310 "Straight Waveguide" sch_x=217 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15156 N$30311 N$30312 "Straight Waveguide" sch_x=217 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15157 N$30313 N$30314 "Straight Waveguide" sch_x=217 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15158 N$30315 N$30316 "Straight Waveguide" sch_x=217 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15159 N$30317 N$30318 "Straight Waveguide" sch_x=217 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15160 N$30319 N$30320 "Straight Waveguide" sch_x=217 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15161 N$30321 N$30322 "Straight Waveguide" sch_x=217 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15162 N$30323 N$30324 "Straight Waveguide" sch_x=217 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15163 N$30325 N$30326 "Straight Waveguide" sch_x=217 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15164 N$30327 N$30328 "Straight Waveguide" sch_x=217 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15165 N$30329 N$30330 "Straight Waveguide" sch_x=217 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15166 N$30331 N$30332 "Straight Waveguide" sch_x=217 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15167 N$30333 N$30334 "Straight Waveguide" sch_x=217 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15168 N$30335 N$30336 "Straight Waveguide" sch_x=217 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15169 N$30337 N$30338 "Straight Waveguide" sch_x=217 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15170 N$30339 N$30340 "Straight Waveguide" sch_x=217 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15171 N$30341 N$30342 "Straight Waveguide" sch_x=217 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15172 N$30343 N$30344 "Straight Waveguide" sch_x=217 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15173 N$30345 N$30346 "Straight Waveguide" sch_x=215 sch_y=43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15174 N$30347 N$30348 "Straight Waveguide" sch_x=215 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15175 N$30349 N$30350 "Straight Waveguide" sch_x=215 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15176 N$30351 N$30352 "Straight Waveguide" sch_x=215 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15177 N$30353 N$30354 "Straight Waveguide" sch_x=215 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15178 N$30355 N$30356 "Straight Waveguide" sch_x=215 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15179 N$30357 N$30358 "Straight Waveguide" sch_x=215 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15180 N$30359 N$30360 "Straight Waveguide" sch_x=215 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15181 N$30361 N$30362 "Straight Waveguide" sch_x=215 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15182 N$30363 N$30364 "Straight Waveguide" sch_x=215 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15183 N$30365 N$30366 "Straight Waveguide" sch_x=215 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15184 N$30367 N$30368 "Straight Waveguide" sch_x=215 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15185 N$30369 N$30370 "Straight Waveguide" sch_x=215 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15186 N$30371 N$30372 "Straight Waveguide" sch_x=215 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15187 N$30373 N$30374 "Straight Waveguide" sch_x=215 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15188 N$30375 N$30376 "Straight Waveguide" sch_x=215 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15189 N$30377 N$30378 "Straight Waveguide" sch_x=215 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15190 N$30379 N$30380 "Straight Waveguide" sch_x=215 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15191 N$30381 N$30382 "Straight Waveguide" sch_x=215 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15192 N$30383 N$30384 "Straight Waveguide" sch_x=215 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15193 N$30385 N$30386 "Straight Waveguide" sch_x=215 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15194 N$30387 N$30388 "Straight Waveguide" sch_x=215 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15195 N$30389 N$30390 "Straight Waveguide" sch_x=215 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15196 N$30391 N$30392 "Straight Waveguide" sch_x=215 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15197 N$30393 N$30394 "Straight Waveguide" sch_x=215 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15198 N$30395 N$30396 "Straight Waveguide" sch_x=215 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15199 N$30397 N$30398 "Straight Waveguide" sch_x=215 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15200 N$30399 N$30400 "Straight Waveguide" sch_x=215 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15201 N$30401 N$30402 "Straight Waveguide" sch_x=215 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15202 N$30403 N$30404 "Straight Waveguide" sch_x=215 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15203 N$30405 N$30406 "Straight Waveguide" sch_x=215 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15204 N$30407 N$30408 "Straight Waveguide" sch_x=215 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15205 N$30409 N$30410 "Straight Waveguide" sch_x=215 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15206 N$30411 N$30412 "Straight Waveguide" sch_x=215 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15207 N$30413 N$30414 "Straight Waveguide" sch_x=215 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15208 N$30415 N$30416 "Straight Waveguide" sch_x=215 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15209 N$30417 N$30418 "Straight Waveguide" sch_x=215 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15210 N$30419 N$30420 "Straight Waveguide" sch_x=215 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15211 N$30421 N$30422 "Straight Waveguide" sch_x=215 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15212 N$30423 N$30424 "Straight Waveguide" sch_x=215 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15213 N$30425 N$30426 "Straight Waveguide" sch_x=215 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15214 N$30427 N$30428 "Straight Waveguide" sch_x=215 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15215 N$30429 N$30430 "Straight Waveguide" sch_x=215 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15216 N$30431 N$30432 "Straight Waveguide" sch_x=215 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15217 N$30433 N$30434 "Straight Waveguide" sch_x=215 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15218 N$30435 N$30436 "Straight Waveguide" sch_x=215 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15219 N$30437 N$30438 "Straight Waveguide" sch_x=215 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15220 N$30439 N$30440 "Straight Waveguide" sch_x=215 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15221 N$30441 N$30442 "Straight Waveguide" sch_x=215 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15222 N$30443 N$30444 "Straight Waveguide" sch_x=215 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15223 N$30445 N$30446 "Straight Waveguide" sch_x=215 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15224 N$30447 N$30448 "Straight Waveguide" sch_x=215 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15225 N$30449 N$30450 "Straight Waveguide" sch_x=215 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15226 N$30451 N$30452 "Straight Waveguide" sch_x=215 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15227 N$30453 N$30454 "Straight Waveguide" sch_x=215 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15228 N$30455 N$30456 "Straight Waveguide" sch_x=215 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15229 N$30457 N$30458 "Straight Waveguide" sch_x=215 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15230 N$30459 N$30460 "Straight Waveguide" sch_x=215 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15231 N$30461 N$30462 "Straight Waveguide" sch_x=215 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15232 N$30463 N$30464 "Straight Waveguide" sch_x=215 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15233 N$30465 N$30466 "Straight Waveguide" sch_x=215 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15234 N$30467 N$30468 "Straight Waveguide" sch_x=215 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15235 N$30469 N$30470 "Straight Waveguide" sch_x=215 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15236 N$30471 N$30472 "Straight Waveguide" sch_x=215 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15237 N$30473 N$30474 "Straight Waveguide" sch_x=215 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15238 N$30475 N$30476 "Straight Waveguide" sch_x=215 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15239 N$30477 N$30478 "Straight Waveguide" sch_x=215 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15240 N$30479 N$30480 "Straight Waveguide" sch_x=215 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15241 N$30481 N$30482 "Straight Waveguide" sch_x=215 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15242 N$30483 N$30484 "Straight Waveguide" sch_x=215 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15243 N$30485 N$30486 "Straight Waveguide" sch_x=215 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15244 N$30487 N$30488 "Straight Waveguide" sch_x=215 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15245 N$30489 N$30490 "Straight Waveguide" sch_x=215 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15246 N$30491 N$30492 "Straight Waveguide" sch_x=215 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15247 N$30493 N$30494 "Straight Waveguide" sch_x=215 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15248 N$30495 N$30496 "Straight Waveguide" sch_x=215 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15249 N$30497 N$30498 "Straight Waveguide" sch_x=215 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15250 N$30499 N$30500 "Straight Waveguide" sch_x=215 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15251 N$30501 N$30502 "Straight Waveguide" sch_x=215 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15252 N$30503 N$30504 "Straight Waveguide" sch_x=215 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15253 N$30505 N$30506 "Straight Waveguide" sch_x=215 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15254 N$30507 N$30508 "Straight Waveguide" sch_x=215 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15255 N$30509 N$30510 "Straight Waveguide" sch_x=215 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15256 N$30511 N$30512 "Straight Waveguide" sch_x=215 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15257 N$30513 N$30514 "Straight Waveguide" sch_x=215 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15258 N$30515 N$30516 "Straight Waveguide" sch_x=215 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15259 N$30517 N$30518 "Straight Waveguide" sch_x=215 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15260 N$30519 N$30520 "Straight Waveguide" sch_x=215 sch_y=-43.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15261 N$30521 N$30522 "Straight Waveguide" sch_x=213 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15262 N$30523 N$30524 "Straight Waveguide" sch_x=213 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15263 N$30525 N$30526 "Straight Waveguide" sch_x=213 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15264 N$30527 N$30528 "Straight Waveguide" sch_x=213 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15265 N$30529 N$30530 "Straight Waveguide" sch_x=213 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15266 N$30531 N$30532 "Straight Waveguide" sch_x=213 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15267 N$30533 N$30534 "Straight Waveguide" sch_x=213 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15268 N$30535 N$30536 "Straight Waveguide" sch_x=213 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15269 N$30537 N$30538 "Straight Waveguide" sch_x=213 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15270 N$30539 N$30540 "Straight Waveguide" sch_x=213 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15271 N$30541 N$30542 "Straight Waveguide" sch_x=213 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15272 N$30543 N$30544 "Straight Waveguide" sch_x=213 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15273 N$30545 N$30546 "Straight Waveguide" sch_x=213 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15274 N$30547 N$30548 "Straight Waveguide" sch_x=213 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15275 N$30549 N$30550 "Straight Waveguide" sch_x=213 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15276 N$30551 N$30552 "Straight Waveguide" sch_x=213 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15277 N$30553 N$30554 "Straight Waveguide" sch_x=213 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15278 N$30555 N$30556 "Straight Waveguide" sch_x=213 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15279 N$30557 N$30558 "Straight Waveguide" sch_x=213 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15280 N$30559 N$30560 "Straight Waveguide" sch_x=213 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15281 N$30561 N$30562 "Straight Waveguide" sch_x=213 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15282 N$30563 N$30564 "Straight Waveguide" sch_x=213 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15283 N$30565 N$30566 "Straight Waveguide" sch_x=213 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15284 N$30567 N$30568 "Straight Waveguide" sch_x=213 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15285 N$30569 N$30570 "Straight Waveguide" sch_x=213 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15286 N$30571 N$30572 "Straight Waveguide" sch_x=213 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15287 N$30573 N$30574 "Straight Waveguide" sch_x=213 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15288 N$30575 N$30576 "Straight Waveguide" sch_x=213 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15289 N$30577 N$30578 "Straight Waveguide" sch_x=213 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15290 N$30579 N$30580 "Straight Waveguide" sch_x=213 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15291 N$30581 N$30582 "Straight Waveguide" sch_x=213 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15292 N$30583 N$30584 "Straight Waveguide" sch_x=213 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15293 N$30585 N$30586 "Straight Waveguide" sch_x=213 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15294 N$30587 N$30588 "Straight Waveguide" sch_x=213 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15295 N$30589 N$30590 "Straight Waveguide" sch_x=213 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15296 N$30591 N$30592 "Straight Waveguide" sch_x=213 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15297 N$30593 N$30594 "Straight Waveguide" sch_x=213 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15298 N$30595 N$30596 "Straight Waveguide" sch_x=213 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15299 N$30597 N$30598 "Straight Waveguide" sch_x=213 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15300 N$30599 N$30600 "Straight Waveguide" sch_x=213 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15301 N$30601 N$30602 "Straight Waveguide" sch_x=213 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15302 N$30603 N$30604 "Straight Waveguide" sch_x=213 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15303 N$30605 N$30606 "Straight Waveguide" sch_x=213 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15304 N$30607 N$30608 "Straight Waveguide" sch_x=213 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15305 N$30609 N$30610 "Straight Waveguide" sch_x=213 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15306 N$30611 N$30612 "Straight Waveguide" sch_x=213 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15307 N$30613 N$30614 "Straight Waveguide" sch_x=213 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15308 N$30615 N$30616 "Straight Waveguide" sch_x=213 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15309 N$30617 N$30618 "Straight Waveguide" sch_x=213 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15310 N$30619 N$30620 "Straight Waveguide" sch_x=213 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15311 N$30621 N$30622 "Straight Waveguide" sch_x=213 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15312 N$30623 N$30624 "Straight Waveguide" sch_x=213 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15313 N$30625 N$30626 "Straight Waveguide" sch_x=213 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15314 N$30627 N$30628 "Straight Waveguide" sch_x=213 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15315 N$30629 N$30630 "Straight Waveguide" sch_x=213 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15316 N$30631 N$30632 "Straight Waveguide" sch_x=213 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15317 N$30633 N$30634 "Straight Waveguide" sch_x=213 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15318 N$30635 N$30636 "Straight Waveguide" sch_x=213 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15319 N$30637 N$30638 "Straight Waveguide" sch_x=213 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15320 N$30639 N$30640 "Straight Waveguide" sch_x=213 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15321 N$30641 N$30642 "Straight Waveguide" sch_x=213 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15322 N$30643 N$30644 "Straight Waveguide" sch_x=213 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15323 N$30645 N$30646 "Straight Waveguide" sch_x=213 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15324 N$30647 N$30648 "Straight Waveguide" sch_x=213 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15325 N$30649 N$30650 "Straight Waveguide" sch_x=213 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15326 N$30651 N$30652 "Straight Waveguide" sch_x=213 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15327 N$30653 N$30654 "Straight Waveguide" sch_x=213 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15328 N$30655 N$30656 "Straight Waveguide" sch_x=213 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15329 N$30657 N$30658 "Straight Waveguide" sch_x=213 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15330 N$30659 N$30660 "Straight Waveguide" sch_x=213 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15331 N$30661 N$30662 "Straight Waveguide" sch_x=213 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15332 N$30663 N$30664 "Straight Waveguide" sch_x=213 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15333 N$30665 N$30666 "Straight Waveguide" sch_x=213 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15334 N$30667 N$30668 "Straight Waveguide" sch_x=213 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15335 N$30669 N$30670 "Straight Waveguide" sch_x=213 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15336 N$30671 N$30672 "Straight Waveguide" sch_x=213 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15337 N$30673 N$30674 "Straight Waveguide" sch_x=213 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15338 N$30675 N$30676 "Straight Waveguide" sch_x=213 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15339 N$30677 N$30678 "Straight Waveguide" sch_x=213 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15340 N$30679 N$30680 "Straight Waveguide" sch_x=213 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15341 N$30681 N$30682 "Straight Waveguide" sch_x=213 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15342 N$30683 N$30684 "Straight Waveguide" sch_x=213 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15343 N$30685 N$30686 "Straight Waveguide" sch_x=213 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15344 N$30687 N$30688 "Straight Waveguide" sch_x=213 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15345 N$30689 N$30690 "Straight Waveguide" sch_x=213 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15346 N$30691 N$30692 "Straight Waveguide" sch_x=213 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15347 N$30693 N$30694 "Straight Waveguide" sch_x=211 sch_y=41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15348 N$30695 N$30696 "Straight Waveguide" sch_x=211 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15349 N$30697 N$30698 "Straight Waveguide" sch_x=211 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15350 N$30699 N$30700 "Straight Waveguide" sch_x=211 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15351 N$30701 N$30702 "Straight Waveguide" sch_x=211 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15352 N$30703 N$30704 "Straight Waveguide" sch_x=211 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15353 N$30705 N$30706 "Straight Waveguide" sch_x=211 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15354 N$30707 N$30708 "Straight Waveguide" sch_x=211 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15355 N$30709 N$30710 "Straight Waveguide" sch_x=211 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15356 N$30711 N$30712 "Straight Waveguide" sch_x=211 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15357 N$30713 N$30714 "Straight Waveguide" sch_x=211 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15358 N$30715 N$30716 "Straight Waveguide" sch_x=211 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15359 N$30717 N$30718 "Straight Waveguide" sch_x=211 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15360 N$30719 N$30720 "Straight Waveguide" sch_x=211 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15361 N$30721 N$30722 "Straight Waveguide" sch_x=211 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15362 N$30723 N$30724 "Straight Waveguide" sch_x=211 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15363 N$30725 N$30726 "Straight Waveguide" sch_x=211 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15364 N$30727 N$30728 "Straight Waveguide" sch_x=211 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15365 N$30729 N$30730 "Straight Waveguide" sch_x=211 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15366 N$30731 N$30732 "Straight Waveguide" sch_x=211 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15367 N$30733 N$30734 "Straight Waveguide" sch_x=211 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15368 N$30735 N$30736 "Straight Waveguide" sch_x=211 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15369 N$30737 N$30738 "Straight Waveguide" sch_x=211 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15370 N$30739 N$30740 "Straight Waveguide" sch_x=211 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15371 N$30741 N$30742 "Straight Waveguide" sch_x=211 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15372 N$30743 N$30744 "Straight Waveguide" sch_x=211 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15373 N$30745 N$30746 "Straight Waveguide" sch_x=211 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15374 N$30747 N$30748 "Straight Waveguide" sch_x=211 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15375 N$30749 N$30750 "Straight Waveguide" sch_x=211 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15376 N$30751 N$30752 "Straight Waveguide" sch_x=211 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15377 N$30753 N$30754 "Straight Waveguide" sch_x=211 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15378 N$30755 N$30756 "Straight Waveguide" sch_x=211 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15379 N$30757 N$30758 "Straight Waveguide" sch_x=211 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15380 N$30759 N$30760 "Straight Waveguide" sch_x=211 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15381 N$30761 N$30762 "Straight Waveguide" sch_x=211 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15382 N$30763 N$30764 "Straight Waveguide" sch_x=211 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15383 N$30765 N$30766 "Straight Waveguide" sch_x=211 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15384 N$30767 N$30768 "Straight Waveguide" sch_x=211 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15385 N$30769 N$30770 "Straight Waveguide" sch_x=211 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15386 N$30771 N$30772 "Straight Waveguide" sch_x=211 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15387 N$30773 N$30774 "Straight Waveguide" sch_x=211 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15388 N$30775 N$30776 "Straight Waveguide" sch_x=211 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15389 N$30777 N$30778 "Straight Waveguide" sch_x=211 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15390 N$30779 N$30780 "Straight Waveguide" sch_x=211 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15391 N$30781 N$30782 "Straight Waveguide" sch_x=211 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15392 N$30783 N$30784 "Straight Waveguide" sch_x=211 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15393 N$30785 N$30786 "Straight Waveguide" sch_x=211 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15394 N$30787 N$30788 "Straight Waveguide" sch_x=211 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15395 N$30789 N$30790 "Straight Waveguide" sch_x=211 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15396 N$30791 N$30792 "Straight Waveguide" sch_x=211 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15397 N$30793 N$30794 "Straight Waveguide" sch_x=211 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15398 N$30795 N$30796 "Straight Waveguide" sch_x=211 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15399 N$30797 N$30798 "Straight Waveguide" sch_x=211 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15400 N$30799 N$30800 "Straight Waveguide" sch_x=211 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15401 N$30801 N$30802 "Straight Waveguide" sch_x=211 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15402 N$30803 N$30804 "Straight Waveguide" sch_x=211 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15403 N$30805 N$30806 "Straight Waveguide" sch_x=211 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15404 N$30807 N$30808 "Straight Waveguide" sch_x=211 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15405 N$30809 N$30810 "Straight Waveguide" sch_x=211 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15406 N$30811 N$30812 "Straight Waveguide" sch_x=211 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15407 N$30813 N$30814 "Straight Waveguide" sch_x=211 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15408 N$30815 N$30816 "Straight Waveguide" sch_x=211 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15409 N$30817 N$30818 "Straight Waveguide" sch_x=211 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15410 N$30819 N$30820 "Straight Waveguide" sch_x=211 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15411 N$30821 N$30822 "Straight Waveguide" sch_x=211 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15412 N$30823 N$30824 "Straight Waveguide" sch_x=211 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15413 N$30825 N$30826 "Straight Waveguide" sch_x=211 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15414 N$30827 N$30828 "Straight Waveguide" sch_x=211 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15415 N$30829 N$30830 "Straight Waveguide" sch_x=211 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15416 N$30831 N$30832 "Straight Waveguide" sch_x=211 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15417 N$30833 N$30834 "Straight Waveguide" sch_x=211 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15418 N$30835 N$30836 "Straight Waveguide" sch_x=211 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15419 N$30837 N$30838 "Straight Waveguide" sch_x=211 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15420 N$30839 N$30840 "Straight Waveguide" sch_x=211 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15421 N$30841 N$30842 "Straight Waveguide" sch_x=211 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15422 N$30843 N$30844 "Straight Waveguide" sch_x=211 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15423 N$30845 N$30846 "Straight Waveguide" sch_x=211 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15424 N$30847 N$30848 "Straight Waveguide" sch_x=211 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15425 N$30849 N$30850 "Straight Waveguide" sch_x=211 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15426 N$30851 N$30852 "Straight Waveguide" sch_x=211 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15427 N$30853 N$30854 "Straight Waveguide" sch_x=211 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15428 N$30855 N$30856 "Straight Waveguide" sch_x=211 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15429 N$30857 N$30858 "Straight Waveguide" sch_x=211 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15430 N$30859 N$30860 "Straight Waveguide" sch_x=211 sch_y=-41.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15431 N$30861 N$30862 "Straight Waveguide" sch_x=209 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15432 N$30863 N$30864 "Straight Waveguide" sch_x=209 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15433 N$30865 N$30866 "Straight Waveguide" sch_x=209 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15434 N$30867 N$30868 "Straight Waveguide" sch_x=209 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15435 N$30869 N$30870 "Straight Waveguide" sch_x=209 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15436 N$30871 N$30872 "Straight Waveguide" sch_x=209 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15437 N$30873 N$30874 "Straight Waveguide" sch_x=209 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15438 N$30875 N$30876 "Straight Waveguide" sch_x=209 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15439 N$30877 N$30878 "Straight Waveguide" sch_x=209 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15440 N$30879 N$30880 "Straight Waveguide" sch_x=209 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15441 N$30881 N$30882 "Straight Waveguide" sch_x=209 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15442 N$30883 N$30884 "Straight Waveguide" sch_x=209 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15443 N$30885 N$30886 "Straight Waveguide" sch_x=209 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15444 N$30887 N$30888 "Straight Waveguide" sch_x=209 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15445 N$30889 N$30890 "Straight Waveguide" sch_x=209 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15446 N$30891 N$30892 "Straight Waveguide" sch_x=209 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15447 N$30893 N$30894 "Straight Waveguide" sch_x=209 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15448 N$30895 N$30896 "Straight Waveguide" sch_x=209 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15449 N$30897 N$30898 "Straight Waveguide" sch_x=209 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15450 N$30899 N$30900 "Straight Waveguide" sch_x=209 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15451 N$30901 N$30902 "Straight Waveguide" sch_x=209 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15452 N$30903 N$30904 "Straight Waveguide" sch_x=209 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15453 N$30905 N$30906 "Straight Waveguide" sch_x=209 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15454 N$30907 N$30908 "Straight Waveguide" sch_x=209 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15455 N$30909 N$30910 "Straight Waveguide" sch_x=209 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15456 N$30911 N$30912 "Straight Waveguide" sch_x=209 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15457 N$30913 N$30914 "Straight Waveguide" sch_x=209 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15458 N$30915 N$30916 "Straight Waveguide" sch_x=209 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15459 N$30917 N$30918 "Straight Waveguide" sch_x=209 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15460 N$30919 N$30920 "Straight Waveguide" sch_x=209 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15461 N$30921 N$30922 "Straight Waveguide" sch_x=209 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15462 N$30923 N$30924 "Straight Waveguide" sch_x=209 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15463 N$30925 N$30926 "Straight Waveguide" sch_x=209 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15464 N$30927 N$30928 "Straight Waveguide" sch_x=209 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15465 N$30929 N$30930 "Straight Waveguide" sch_x=209 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15466 N$30931 N$30932 "Straight Waveguide" sch_x=209 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15467 N$30933 N$30934 "Straight Waveguide" sch_x=209 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15468 N$30935 N$30936 "Straight Waveguide" sch_x=209 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15469 N$30937 N$30938 "Straight Waveguide" sch_x=209 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15470 N$30939 N$30940 "Straight Waveguide" sch_x=209 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15471 N$30941 N$30942 "Straight Waveguide" sch_x=209 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15472 N$30943 N$30944 "Straight Waveguide" sch_x=209 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15473 N$30945 N$30946 "Straight Waveguide" sch_x=209 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15474 N$30947 N$30948 "Straight Waveguide" sch_x=209 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15475 N$30949 N$30950 "Straight Waveguide" sch_x=209 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15476 N$30951 N$30952 "Straight Waveguide" sch_x=209 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15477 N$30953 N$30954 "Straight Waveguide" sch_x=209 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15478 N$30955 N$30956 "Straight Waveguide" sch_x=209 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15479 N$30957 N$30958 "Straight Waveguide" sch_x=209 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15480 N$30959 N$30960 "Straight Waveguide" sch_x=209 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15481 N$30961 N$30962 "Straight Waveguide" sch_x=209 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15482 N$30963 N$30964 "Straight Waveguide" sch_x=209 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15483 N$30965 N$30966 "Straight Waveguide" sch_x=209 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15484 N$30967 N$30968 "Straight Waveguide" sch_x=209 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15485 N$30969 N$30970 "Straight Waveguide" sch_x=209 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15486 N$30971 N$30972 "Straight Waveguide" sch_x=209 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15487 N$30973 N$30974 "Straight Waveguide" sch_x=209 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15488 N$30975 N$30976 "Straight Waveguide" sch_x=209 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15489 N$30977 N$30978 "Straight Waveguide" sch_x=209 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15490 N$30979 N$30980 "Straight Waveguide" sch_x=209 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15491 N$30981 N$30982 "Straight Waveguide" sch_x=209 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15492 N$30983 N$30984 "Straight Waveguide" sch_x=209 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15493 N$30985 N$30986 "Straight Waveguide" sch_x=209 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15494 N$30987 N$30988 "Straight Waveguide" sch_x=209 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15495 N$30989 N$30990 "Straight Waveguide" sch_x=209 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15496 N$30991 N$30992 "Straight Waveguide" sch_x=209 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15497 N$30993 N$30994 "Straight Waveguide" sch_x=209 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15498 N$30995 N$30996 "Straight Waveguide" sch_x=209 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15499 N$30997 N$30998 "Straight Waveguide" sch_x=209 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15500 N$30999 N$31000 "Straight Waveguide" sch_x=209 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15501 N$31001 N$31002 "Straight Waveguide" sch_x=209 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15502 N$31003 N$31004 "Straight Waveguide" sch_x=209 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15503 N$31005 N$31006 "Straight Waveguide" sch_x=209 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15504 N$31007 N$31008 "Straight Waveguide" sch_x=209 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15505 N$31009 N$31010 "Straight Waveguide" sch_x=209 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15506 N$31011 N$31012 "Straight Waveguide" sch_x=209 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15507 N$31013 N$31014 "Straight Waveguide" sch_x=209 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15508 N$31015 N$31016 "Straight Waveguide" sch_x=209 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15509 N$31017 N$31018 "Straight Waveguide" sch_x=209 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15510 N$31019 N$31020 "Straight Waveguide" sch_x=209 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15511 N$31021 N$31022 "Straight Waveguide" sch_x=209 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15512 N$31023 N$31024 "Straight Waveguide" sch_x=209 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15513 N$31025 N$31026 "Straight Waveguide" sch_x=207 sch_y=39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15514 N$31027 N$31028 "Straight Waveguide" sch_x=207 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15515 N$31029 N$31030 "Straight Waveguide" sch_x=207 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15516 N$31031 N$31032 "Straight Waveguide" sch_x=207 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15517 N$31033 N$31034 "Straight Waveguide" sch_x=207 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15518 N$31035 N$31036 "Straight Waveguide" sch_x=207 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15519 N$31037 N$31038 "Straight Waveguide" sch_x=207 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15520 N$31039 N$31040 "Straight Waveguide" sch_x=207 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15521 N$31041 N$31042 "Straight Waveguide" sch_x=207 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15522 N$31043 N$31044 "Straight Waveguide" sch_x=207 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15523 N$31045 N$31046 "Straight Waveguide" sch_x=207 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15524 N$31047 N$31048 "Straight Waveguide" sch_x=207 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15525 N$31049 N$31050 "Straight Waveguide" sch_x=207 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15526 N$31051 N$31052 "Straight Waveguide" sch_x=207 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15527 N$31053 N$31054 "Straight Waveguide" sch_x=207 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15528 N$31055 N$31056 "Straight Waveguide" sch_x=207 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15529 N$31057 N$31058 "Straight Waveguide" sch_x=207 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15530 N$31059 N$31060 "Straight Waveguide" sch_x=207 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15531 N$31061 N$31062 "Straight Waveguide" sch_x=207 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15532 N$31063 N$31064 "Straight Waveguide" sch_x=207 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15533 N$31065 N$31066 "Straight Waveguide" sch_x=207 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15534 N$31067 N$31068 "Straight Waveguide" sch_x=207 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15535 N$31069 N$31070 "Straight Waveguide" sch_x=207 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15536 N$31071 N$31072 "Straight Waveguide" sch_x=207 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15537 N$31073 N$31074 "Straight Waveguide" sch_x=207 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15538 N$31075 N$31076 "Straight Waveguide" sch_x=207 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15539 N$31077 N$31078 "Straight Waveguide" sch_x=207 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15540 N$31079 N$31080 "Straight Waveguide" sch_x=207 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15541 N$31081 N$31082 "Straight Waveguide" sch_x=207 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15542 N$31083 N$31084 "Straight Waveguide" sch_x=207 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15543 N$31085 N$31086 "Straight Waveguide" sch_x=207 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15544 N$31087 N$31088 "Straight Waveguide" sch_x=207 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15545 N$31089 N$31090 "Straight Waveguide" sch_x=207 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15546 N$31091 N$31092 "Straight Waveguide" sch_x=207 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15547 N$31093 N$31094 "Straight Waveguide" sch_x=207 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15548 N$31095 N$31096 "Straight Waveguide" sch_x=207 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15549 N$31097 N$31098 "Straight Waveguide" sch_x=207 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15550 N$31099 N$31100 "Straight Waveguide" sch_x=207 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15551 N$31101 N$31102 "Straight Waveguide" sch_x=207 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15552 N$31103 N$31104 "Straight Waveguide" sch_x=207 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15553 N$31105 N$31106 "Straight Waveguide" sch_x=207 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15554 N$31107 N$31108 "Straight Waveguide" sch_x=207 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15555 N$31109 N$31110 "Straight Waveguide" sch_x=207 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15556 N$31111 N$31112 "Straight Waveguide" sch_x=207 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15557 N$31113 N$31114 "Straight Waveguide" sch_x=207 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15558 N$31115 N$31116 "Straight Waveguide" sch_x=207 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15559 N$31117 N$31118 "Straight Waveguide" sch_x=207 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15560 N$31119 N$31120 "Straight Waveguide" sch_x=207 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15561 N$31121 N$31122 "Straight Waveguide" sch_x=207 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15562 N$31123 N$31124 "Straight Waveguide" sch_x=207 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15563 N$31125 N$31126 "Straight Waveguide" sch_x=207 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15564 N$31127 N$31128 "Straight Waveguide" sch_x=207 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15565 N$31129 N$31130 "Straight Waveguide" sch_x=207 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15566 N$31131 N$31132 "Straight Waveguide" sch_x=207 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15567 N$31133 N$31134 "Straight Waveguide" sch_x=207 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15568 N$31135 N$31136 "Straight Waveguide" sch_x=207 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15569 N$31137 N$31138 "Straight Waveguide" sch_x=207 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15570 N$31139 N$31140 "Straight Waveguide" sch_x=207 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15571 N$31141 N$31142 "Straight Waveguide" sch_x=207 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15572 N$31143 N$31144 "Straight Waveguide" sch_x=207 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15573 N$31145 N$31146 "Straight Waveguide" sch_x=207 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15574 N$31147 N$31148 "Straight Waveguide" sch_x=207 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15575 N$31149 N$31150 "Straight Waveguide" sch_x=207 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15576 N$31151 N$31152 "Straight Waveguide" sch_x=207 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15577 N$31153 N$31154 "Straight Waveguide" sch_x=207 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15578 N$31155 N$31156 "Straight Waveguide" sch_x=207 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15579 N$31157 N$31158 "Straight Waveguide" sch_x=207 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15580 N$31159 N$31160 "Straight Waveguide" sch_x=207 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15581 N$31161 N$31162 "Straight Waveguide" sch_x=207 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15582 N$31163 N$31164 "Straight Waveguide" sch_x=207 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15583 N$31165 N$31166 "Straight Waveguide" sch_x=207 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15584 N$31167 N$31168 "Straight Waveguide" sch_x=207 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15585 N$31169 N$31170 "Straight Waveguide" sch_x=207 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15586 N$31171 N$31172 "Straight Waveguide" sch_x=207 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15587 N$31173 N$31174 "Straight Waveguide" sch_x=207 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15588 N$31175 N$31176 "Straight Waveguide" sch_x=207 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15589 N$31177 N$31178 "Straight Waveguide" sch_x=207 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15590 N$31179 N$31180 "Straight Waveguide" sch_x=207 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15591 N$31181 N$31182 "Straight Waveguide" sch_x=207 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15592 N$31183 N$31184 "Straight Waveguide" sch_x=207 sch_y=-39.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15593 N$31185 N$31186 "Straight Waveguide" sch_x=205 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15594 N$31187 N$31188 "Straight Waveguide" sch_x=205 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15595 N$31189 N$31190 "Straight Waveguide" sch_x=205 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15596 N$31191 N$31192 "Straight Waveguide" sch_x=205 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15597 N$31193 N$31194 "Straight Waveguide" sch_x=205 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15598 N$31195 N$31196 "Straight Waveguide" sch_x=205 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15599 N$31197 N$31198 "Straight Waveguide" sch_x=205 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15600 N$31199 N$31200 "Straight Waveguide" sch_x=205 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15601 N$31201 N$31202 "Straight Waveguide" sch_x=205 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15602 N$31203 N$31204 "Straight Waveguide" sch_x=205 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15603 N$31205 N$31206 "Straight Waveguide" sch_x=205 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15604 N$31207 N$31208 "Straight Waveguide" sch_x=205 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15605 N$31209 N$31210 "Straight Waveguide" sch_x=205 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15606 N$31211 N$31212 "Straight Waveguide" sch_x=205 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15607 N$31213 N$31214 "Straight Waveguide" sch_x=205 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15608 N$31215 N$31216 "Straight Waveguide" sch_x=205 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15609 N$31217 N$31218 "Straight Waveguide" sch_x=205 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15610 N$31219 N$31220 "Straight Waveguide" sch_x=205 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15611 N$31221 N$31222 "Straight Waveguide" sch_x=205 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15612 N$31223 N$31224 "Straight Waveguide" sch_x=205 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15613 N$31225 N$31226 "Straight Waveguide" sch_x=205 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15614 N$31227 N$31228 "Straight Waveguide" sch_x=205 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15615 N$31229 N$31230 "Straight Waveguide" sch_x=205 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15616 N$31231 N$31232 "Straight Waveguide" sch_x=205 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15617 N$31233 N$31234 "Straight Waveguide" sch_x=205 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15618 N$31235 N$31236 "Straight Waveguide" sch_x=205 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15619 N$31237 N$31238 "Straight Waveguide" sch_x=205 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15620 N$31239 N$31240 "Straight Waveguide" sch_x=205 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15621 N$31241 N$31242 "Straight Waveguide" sch_x=205 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15622 N$31243 N$31244 "Straight Waveguide" sch_x=205 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15623 N$31245 N$31246 "Straight Waveguide" sch_x=205 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15624 N$31247 N$31248 "Straight Waveguide" sch_x=205 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15625 N$31249 N$31250 "Straight Waveguide" sch_x=205 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15626 N$31251 N$31252 "Straight Waveguide" sch_x=205 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15627 N$31253 N$31254 "Straight Waveguide" sch_x=205 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15628 N$31255 N$31256 "Straight Waveguide" sch_x=205 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15629 N$31257 N$31258 "Straight Waveguide" sch_x=205 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15630 N$31259 N$31260 "Straight Waveguide" sch_x=205 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15631 N$31261 N$31262 "Straight Waveguide" sch_x=205 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15632 N$31263 N$31264 "Straight Waveguide" sch_x=205 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15633 N$31265 N$31266 "Straight Waveguide" sch_x=205 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15634 N$31267 N$31268 "Straight Waveguide" sch_x=205 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15635 N$31269 N$31270 "Straight Waveguide" sch_x=205 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15636 N$31271 N$31272 "Straight Waveguide" sch_x=205 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15637 N$31273 N$31274 "Straight Waveguide" sch_x=205 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15638 N$31275 N$31276 "Straight Waveguide" sch_x=205 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15639 N$31277 N$31278 "Straight Waveguide" sch_x=205 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15640 N$31279 N$31280 "Straight Waveguide" sch_x=205 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15641 N$31281 N$31282 "Straight Waveguide" sch_x=205 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15642 N$31283 N$31284 "Straight Waveguide" sch_x=205 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15643 N$31285 N$31286 "Straight Waveguide" sch_x=205 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15644 N$31287 N$31288 "Straight Waveguide" sch_x=205 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15645 N$31289 N$31290 "Straight Waveguide" sch_x=205 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15646 N$31291 N$31292 "Straight Waveguide" sch_x=205 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15647 N$31293 N$31294 "Straight Waveguide" sch_x=205 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15648 N$31295 N$31296 "Straight Waveguide" sch_x=205 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15649 N$31297 N$31298 "Straight Waveguide" sch_x=205 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15650 N$31299 N$31300 "Straight Waveguide" sch_x=205 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15651 N$31301 N$31302 "Straight Waveguide" sch_x=205 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15652 N$31303 N$31304 "Straight Waveguide" sch_x=205 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15653 N$31305 N$31306 "Straight Waveguide" sch_x=205 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15654 N$31307 N$31308 "Straight Waveguide" sch_x=205 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15655 N$31309 N$31310 "Straight Waveguide" sch_x=205 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15656 N$31311 N$31312 "Straight Waveguide" sch_x=205 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15657 N$31313 N$31314 "Straight Waveguide" sch_x=205 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15658 N$31315 N$31316 "Straight Waveguide" sch_x=205 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15659 N$31317 N$31318 "Straight Waveguide" sch_x=205 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15660 N$31319 N$31320 "Straight Waveguide" sch_x=205 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15661 N$31321 N$31322 "Straight Waveguide" sch_x=205 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15662 N$31323 N$31324 "Straight Waveguide" sch_x=205 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15663 N$31325 N$31326 "Straight Waveguide" sch_x=205 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15664 N$31327 N$31328 "Straight Waveguide" sch_x=205 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15665 N$31329 N$31330 "Straight Waveguide" sch_x=205 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15666 N$31331 N$31332 "Straight Waveguide" sch_x=205 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15667 N$31333 N$31334 "Straight Waveguide" sch_x=205 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15668 N$31335 N$31336 "Straight Waveguide" sch_x=205 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15669 N$31337 N$31338 "Straight Waveguide" sch_x=205 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15670 N$31339 N$31340 "Straight Waveguide" sch_x=205 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15671 N$31341 N$31342 "Straight Waveguide" sch_x=203 sch_y=37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15672 N$31343 N$31344 "Straight Waveguide" sch_x=203 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15673 N$31345 N$31346 "Straight Waveguide" sch_x=203 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15674 N$31347 N$31348 "Straight Waveguide" sch_x=203 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15675 N$31349 N$31350 "Straight Waveguide" sch_x=203 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15676 N$31351 N$31352 "Straight Waveguide" sch_x=203 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15677 N$31353 N$31354 "Straight Waveguide" sch_x=203 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15678 N$31355 N$31356 "Straight Waveguide" sch_x=203 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15679 N$31357 N$31358 "Straight Waveguide" sch_x=203 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15680 N$31359 N$31360 "Straight Waveguide" sch_x=203 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15681 N$31361 N$31362 "Straight Waveguide" sch_x=203 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15682 N$31363 N$31364 "Straight Waveguide" sch_x=203 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15683 N$31365 N$31366 "Straight Waveguide" sch_x=203 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15684 N$31367 N$31368 "Straight Waveguide" sch_x=203 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15685 N$31369 N$31370 "Straight Waveguide" sch_x=203 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15686 N$31371 N$31372 "Straight Waveguide" sch_x=203 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15687 N$31373 N$31374 "Straight Waveguide" sch_x=203 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15688 N$31375 N$31376 "Straight Waveguide" sch_x=203 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15689 N$31377 N$31378 "Straight Waveguide" sch_x=203 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15690 N$31379 N$31380 "Straight Waveguide" sch_x=203 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15691 N$31381 N$31382 "Straight Waveguide" sch_x=203 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15692 N$31383 N$31384 "Straight Waveguide" sch_x=203 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15693 N$31385 N$31386 "Straight Waveguide" sch_x=203 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15694 N$31387 N$31388 "Straight Waveguide" sch_x=203 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15695 N$31389 N$31390 "Straight Waveguide" sch_x=203 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15696 N$31391 N$31392 "Straight Waveguide" sch_x=203 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15697 N$31393 N$31394 "Straight Waveguide" sch_x=203 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15698 N$31395 N$31396 "Straight Waveguide" sch_x=203 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15699 N$31397 N$31398 "Straight Waveguide" sch_x=203 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15700 N$31399 N$31400 "Straight Waveguide" sch_x=203 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15701 N$31401 N$31402 "Straight Waveguide" sch_x=203 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15702 N$31403 N$31404 "Straight Waveguide" sch_x=203 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15703 N$31405 N$31406 "Straight Waveguide" sch_x=203 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15704 N$31407 N$31408 "Straight Waveguide" sch_x=203 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15705 N$31409 N$31410 "Straight Waveguide" sch_x=203 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15706 N$31411 N$31412 "Straight Waveguide" sch_x=203 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15707 N$31413 N$31414 "Straight Waveguide" sch_x=203 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15708 N$31415 N$31416 "Straight Waveguide" sch_x=203 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15709 N$31417 N$31418 "Straight Waveguide" sch_x=203 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15710 N$31419 N$31420 "Straight Waveguide" sch_x=203 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15711 N$31421 N$31422 "Straight Waveguide" sch_x=203 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15712 N$31423 N$31424 "Straight Waveguide" sch_x=203 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15713 N$31425 N$31426 "Straight Waveguide" sch_x=203 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15714 N$31427 N$31428 "Straight Waveguide" sch_x=203 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15715 N$31429 N$31430 "Straight Waveguide" sch_x=203 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15716 N$31431 N$31432 "Straight Waveguide" sch_x=203 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15717 N$31433 N$31434 "Straight Waveguide" sch_x=203 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15718 N$31435 N$31436 "Straight Waveguide" sch_x=203 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15719 N$31437 N$31438 "Straight Waveguide" sch_x=203 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15720 N$31439 N$31440 "Straight Waveguide" sch_x=203 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15721 N$31441 N$31442 "Straight Waveguide" sch_x=203 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15722 N$31443 N$31444 "Straight Waveguide" sch_x=203 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15723 N$31445 N$31446 "Straight Waveguide" sch_x=203 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15724 N$31447 N$31448 "Straight Waveguide" sch_x=203 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15725 N$31449 N$31450 "Straight Waveguide" sch_x=203 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15726 N$31451 N$31452 "Straight Waveguide" sch_x=203 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15727 N$31453 N$31454 "Straight Waveguide" sch_x=203 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15728 N$31455 N$31456 "Straight Waveguide" sch_x=203 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15729 N$31457 N$31458 "Straight Waveguide" sch_x=203 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15730 N$31459 N$31460 "Straight Waveguide" sch_x=203 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15731 N$31461 N$31462 "Straight Waveguide" sch_x=203 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15732 N$31463 N$31464 "Straight Waveguide" sch_x=203 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15733 N$31465 N$31466 "Straight Waveguide" sch_x=203 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15734 N$31467 N$31468 "Straight Waveguide" sch_x=203 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15735 N$31469 N$31470 "Straight Waveguide" sch_x=203 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15736 N$31471 N$31472 "Straight Waveguide" sch_x=203 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15737 N$31473 N$31474 "Straight Waveguide" sch_x=203 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15738 N$31475 N$31476 "Straight Waveguide" sch_x=203 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15739 N$31477 N$31478 "Straight Waveguide" sch_x=203 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15740 N$31479 N$31480 "Straight Waveguide" sch_x=203 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15741 N$31481 N$31482 "Straight Waveguide" sch_x=203 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15742 N$31483 N$31484 "Straight Waveguide" sch_x=203 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15743 N$31485 N$31486 "Straight Waveguide" sch_x=203 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15744 N$31487 N$31488 "Straight Waveguide" sch_x=203 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15745 N$31489 N$31490 "Straight Waveguide" sch_x=203 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15746 N$31491 N$31492 "Straight Waveguide" sch_x=203 sch_y=-37.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15747 N$31493 N$31494 "Straight Waveguide" sch_x=201 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15748 N$31495 N$31496 "Straight Waveguide" sch_x=201 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15749 N$31497 N$31498 "Straight Waveguide" sch_x=201 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15750 N$31499 N$31500 "Straight Waveguide" sch_x=201 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15751 N$31501 N$31502 "Straight Waveguide" sch_x=201 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15752 N$31503 N$31504 "Straight Waveguide" sch_x=201 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15753 N$31505 N$31506 "Straight Waveguide" sch_x=201 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15754 N$31507 N$31508 "Straight Waveguide" sch_x=201 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15755 N$31509 N$31510 "Straight Waveguide" sch_x=201 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15756 N$31511 N$31512 "Straight Waveguide" sch_x=201 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15757 N$31513 N$31514 "Straight Waveguide" sch_x=201 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15758 N$31515 N$31516 "Straight Waveguide" sch_x=201 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15759 N$31517 N$31518 "Straight Waveguide" sch_x=201 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15760 N$31519 N$31520 "Straight Waveguide" sch_x=201 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15761 N$31521 N$31522 "Straight Waveguide" sch_x=201 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15762 N$31523 N$31524 "Straight Waveguide" sch_x=201 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15763 N$31525 N$31526 "Straight Waveguide" sch_x=201 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15764 N$31527 N$31528 "Straight Waveguide" sch_x=201 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15765 N$31529 N$31530 "Straight Waveguide" sch_x=201 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15766 N$31531 N$31532 "Straight Waveguide" sch_x=201 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15767 N$31533 N$31534 "Straight Waveguide" sch_x=201 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15768 N$31535 N$31536 "Straight Waveguide" sch_x=201 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15769 N$31537 N$31538 "Straight Waveguide" sch_x=201 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15770 N$31539 N$31540 "Straight Waveguide" sch_x=201 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15771 N$31541 N$31542 "Straight Waveguide" sch_x=201 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15772 N$31543 N$31544 "Straight Waveguide" sch_x=201 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15773 N$31545 N$31546 "Straight Waveguide" sch_x=201 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15774 N$31547 N$31548 "Straight Waveguide" sch_x=201 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15775 N$31549 N$31550 "Straight Waveguide" sch_x=201 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15776 N$31551 N$31552 "Straight Waveguide" sch_x=201 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15777 N$31553 N$31554 "Straight Waveguide" sch_x=201 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15778 N$31555 N$31556 "Straight Waveguide" sch_x=201 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15779 N$31557 N$31558 "Straight Waveguide" sch_x=201 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15780 N$31559 N$31560 "Straight Waveguide" sch_x=201 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15781 N$31561 N$31562 "Straight Waveguide" sch_x=201 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15782 N$31563 N$31564 "Straight Waveguide" sch_x=201 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15783 N$31565 N$31566 "Straight Waveguide" sch_x=201 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15784 N$31567 N$31568 "Straight Waveguide" sch_x=201 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15785 N$31569 N$31570 "Straight Waveguide" sch_x=201 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15786 N$31571 N$31572 "Straight Waveguide" sch_x=201 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15787 N$31573 N$31574 "Straight Waveguide" sch_x=201 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15788 N$31575 N$31576 "Straight Waveguide" sch_x=201 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15789 N$31577 N$31578 "Straight Waveguide" sch_x=201 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15790 N$31579 N$31580 "Straight Waveguide" sch_x=201 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15791 N$31581 N$31582 "Straight Waveguide" sch_x=201 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15792 N$31583 N$31584 "Straight Waveguide" sch_x=201 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15793 N$31585 N$31586 "Straight Waveguide" sch_x=201 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15794 N$31587 N$31588 "Straight Waveguide" sch_x=201 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15795 N$31589 N$31590 "Straight Waveguide" sch_x=201 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15796 N$31591 N$31592 "Straight Waveguide" sch_x=201 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15797 N$31593 N$31594 "Straight Waveguide" sch_x=201 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15798 N$31595 N$31596 "Straight Waveguide" sch_x=201 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15799 N$31597 N$31598 "Straight Waveguide" sch_x=201 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15800 N$31599 N$31600 "Straight Waveguide" sch_x=201 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15801 N$31601 N$31602 "Straight Waveguide" sch_x=201 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15802 N$31603 N$31604 "Straight Waveguide" sch_x=201 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15803 N$31605 N$31606 "Straight Waveguide" sch_x=201 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15804 N$31607 N$31608 "Straight Waveguide" sch_x=201 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15805 N$31609 N$31610 "Straight Waveguide" sch_x=201 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15806 N$31611 N$31612 "Straight Waveguide" sch_x=201 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15807 N$31613 N$31614 "Straight Waveguide" sch_x=201 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15808 N$31615 N$31616 "Straight Waveguide" sch_x=201 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15809 N$31617 N$31618 "Straight Waveguide" sch_x=201 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15810 N$31619 N$31620 "Straight Waveguide" sch_x=201 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15811 N$31621 N$31622 "Straight Waveguide" sch_x=201 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15812 N$31623 N$31624 "Straight Waveguide" sch_x=201 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15813 N$31625 N$31626 "Straight Waveguide" sch_x=201 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15814 N$31627 N$31628 "Straight Waveguide" sch_x=201 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15815 N$31629 N$31630 "Straight Waveguide" sch_x=201 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15816 N$31631 N$31632 "Straight Waveguide" sch_x=201 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15817 N$31633 N$31634 "Straight Waveguide" sch_x=201 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15818 N$31635 N$31636 "Straight Waveguide" sch_x=201 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15819 N$31637 N$31638 "Straight Waveguide" sch_x=201 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15820 N$31639 N$31640 "Straight Waveguide" sch_x=201 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15821 N$31641 N$31642 "Straight Waveguide" sch_x=199 sch_y=35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15822 N$31643 N$31644 "Straight Waveguide" sch_x=199 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15823 N$31645 N$31646 "Straight Waveguide" sch_x=199 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15824 N$31647 N$31648 "Straight Waveguide" sch_x=199 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15825 N$31649 N$31650 "Straight Waveguide" sch_x=199 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15826 N$31651 N$31652 "Straight Waveguide" sch_x=199 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15827 N$31653 N$31654 "Straight Waveguide" sch_x=199 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15828 N$31655 N$31656 "Straight Waveguide" sch_x=199 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15829 N$31657 N$31658 "Straight Waveguide" sch_x=199 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15830 N$31659 N$31660 "Straight Waveguide" sch_x=199 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15831 N$31661 N$31662 "Straight Waveguide" sch_x=199 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15832 N$31663 N$31664 "Straight Waveguide" sch_x=199 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15833 N$31665 N$31666 "Straight Waveguide" sch_x=199 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15834 N$31667 N$31668 "Straight Waveguide" sch_x=199 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15835 N$31669 N$31670 "Straight Waveguide" sch_x=199 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15836 N$31671 N$31672 "Straight Waveguide" sch_x=199 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15837 N$31673 N$31674 "Straight Waveguide" sch_x=199 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15838 N$31675 N$31676 "Straight Waveguide" sch_x=199 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15839 N$31677 N$31678 "Straight Waveguide" sch_x=199 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15840 N$31679 N$31680 "Straight Waveguide" sch_x=199 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15841 N$31681 N$31682 "Straight Waveguide" sch_x=199 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15842 N$31683 N$31684 "Straight Waveguide" sch_x=199 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15843 N$31685 N$31686 "Straight Waveguide" sch_x=199 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15844 N$31687 N$31688 "Straight Waveguide" sch_x=199 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15845 N$31689 N$31690 "Straight Waveguide" sch_x=199 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15846 N$31691 N$31692 "Straight Waveguide" sch_x=199 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15847 N$31693 N$31694 "Straight Waveguide" sch_x=199 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15848 N$31695 N$31696 "Straight Waveguide" sch_x=199 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15849 N$31697 N$31698 "Straight Waveguide" sch_x=199 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15850 N$31699 N$31700 "Straight Waveguide" sch_x=199 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15851 N$31701 N$31702 "Straight Waveguide" sch_x=199 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15852 N$31703 N$31704 "Straight Waveguide" sch_x=199 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15853 N$31705 N$31706 "Straight Waveguide" sch_x=199 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15854 N$31707 N$31708 "Straight Waveguide" sch_x=199 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15855 N$31709 N$31710 "Straight Waveguide" sch_x=199 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15856 N$31711 N$31712 "Straight Waveguide" sch_x=199 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15857 N$31713 N$31714 "Straight Waveguide" sch_x=199 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15858 N$31715 N$31716 "Straight Waveguide" sch_x=199 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15859 N$31717 N$31718 "Straight Waveguide" sch_x=199 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15860 N$31719 N$31720 "Straight Waveguide" sch_x=199 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15861 N$31721 N$31722 "Straight Waveguide" sch_x=199 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15862 N$31723 N$31724 "Straight Waveguide" sch_x=199 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15863 N$31725 N$31726 "Straight Waveguide" sch_x=199 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15864 N$31727 N$31728 "Straight Waveguide" sch_x=199 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15865 N$31729 N$31730 "Straight Waveguide" sch_x=199 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15866 N$31731 N$31732 "Straight Waveguide" sch_x=199 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15867 N$31733 N$31734 "Straight Waveguide" sch_x=199 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15868 N$31735 N$31736 "Straight Waveguide" sch_x=199 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15869 N$31737 N$31738 "Straight Waveguide" sch_x=199 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15870 N$31739 N$31740 "Straight Waveguide" sch_x=199 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15871 N$31741 N$31742 "Straight Waveguide" sch_x=199 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15872 N$31743 N$31744 "Straight Waveguide" sch_x=199 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15873 N$31745 N$31746 "Straight Waveguide" sch_x=199 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15874 N$31747 N$31748 "Straight Waveguide" sch_x=199 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15875 N$31749 N$31750 "Straight Waveguide" sch_x=199 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15876 N$31751 N$31752 "Straight Waveguide" sch_x=199 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15877 N$31753 N$31754 "Straight Waveguide" sch_x=199 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15878 N$31755 N$31756 "Straight Waveguide" sch_x=199 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15879 N$31757 N$31758 "Straight Waveguide" sch_x=199 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15880 N$31759 N$31760 "Straight Waveguide" sch_x=199 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15881 N$31761 N$31762 "Straight Waveguide" sch_x=199 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15882 N$31763 N$31764 "Straight Waveguide" sch_x=199 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15883 N$31765 N$31766 "Straight Waveguide" sch_x=199 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15884 N$31767 N$31768 "Straight Waveguide" sch_x=199 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15885 N$31769 N$31770 "Straight Waveguide" sch_x=199 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15886 N$31771 N$31772 "Straight Waveguide" sch_x=199 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15887 N$31773 N$31774 "Straight Waveguide" sch_x=199 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15888 N$31775 N$31776 "Straight Waveguide" sch_x=199 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15889 N$31777 N$31778 "Straight Waveguide" sch_x=199 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15890 N$31779 N$31780 "Straight Waveguide" sch_x=199 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15891 N$31781 N$31782 "Straight Waveguide" sch_x=199 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15892 N$31783 N$31784 "Straight Waveguide" sch_x=199 sch_y=-35.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15893 N$31785 N$31786 "Straight Waveguide" sch_x=197 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15894 N$31787 N$31788 "Straight Waveguide" sch_x=197 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15895 N$31789 N$31790 "Straight Waveguide" sch_x=197 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15896 N$31791 N$31792 "Straight Waveguide" sch_x=197 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15897 N$31793 N$31794 "Straight Waveguide" sch_x=197 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15898 N$31795 N$31796 "Straight Waveguide" sch_x=197 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15899 N$31797 N$31798 "Straight Waveguide" sch_x=197 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15900 N$31799 N$31800 "Straight Waveguide" sch_x=197 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15901 N$31801 N$31802 "Straight Waveguide" sch_x=197 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15902 N$31803 N$31804 "Straight Waveguide" sch_x=197 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15903 N$31805 N$31806 "Straight Waveguide" sch_x=197 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15904 N$31807 N$31808 "Straight Waveguide" sch_x=197 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15905 N$31809 N$31810 "Straight Waveguide" sch_x=197 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15906 N$31811 N$31812 "Straight Waveguide" sch_x=197 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15907 N$31813 N$31814 "Straight Waveguide" sch_x=197 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15908 N$31815 N$31816 "Straight Waveguide" sch_x=197 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15909 N$31817 N$31818 "Straight Waveguide" sch_x=197 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15910 N$31819 N$31820 "Straight Waveguide" sch_x=197 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15911 N$31821 N$31822 "Straight Waveguide" sch_x=197 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15912 N$31823 N$31824 "Straight Waveguide" sch_x=197 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15913 N$31825 N$31826 "Straight Waveguide" sch_x=197 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15914 N$31827 N$31828 "Straight Waveguide" sch_x=197 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15915 N$31829 N$31830 "Straight Waveguide" sch_x=197 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15916 N$31831 N$31832 "Straight Waveguide" sch_x=197 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15917 N$31833 N$31834 "Straight Waveguide" sch_x=197 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15918 N$31835 N$31836 "Straight Waveguide" sch_x=197 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15919 N$31837 N$31838 "Straight Waveguide" sch_x=197 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15920 N$31839 N$31840 "Straight Waveguide" sch_x=197 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15921 N$31841 N$31842 "Straight Waveguide" sch_x=197 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15922 N$31843 N$31844 "Straight Waveguide" sch_x=197 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15923 N$31845 N$31846 "Straight Waveguide" sch_x=197 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15924 N$31847 N$31848 "Straight Waveguide" sch_x=197 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15925 N$31849 N$31850 "Straight Waveguide" sch_x=197 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15926 N$31851 N$31852 "Straight Waveguide" sch_x=197 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15927 N$31853 N$31854 "Straight Waveguide" sch_x=197 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15928 N$31855 N$31856 "Straight Waveguide" sch_x=197 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15929 N$31857 N$31858 "Straight Waveguide" sch_x=197 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15930 N$31859 N$31860 "Straight Waveguide" sch_x=197 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15931 N$31861 N$31862 "Straight Waveguide" sch_x=197 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15932 N$31863 N$31864 "Straight Waveguide" sch_x=197 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15933 N$31865 N$31866 "Straight Waveguide" sch_x=197 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15934 N$31867 N$31868 "Straight Waveguide" sch_x=197 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15935 N$31869 N$31870 "Straight Waveguide" sch_x=197 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15936 N$31871 N$31872 "Straight Waveguide" sch_x=197 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15937 N$31873 N$31874 "Straight Waveguide" sch_x=197 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15938 N$31875 N$31876 "Straight Waveguide" sch_x=197 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15939 N$31877 N$31878 "Straight Waveguide" sch_x=197 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15940 N$31879 N$31880 "Straight Waveguide" sch_x=197 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15941 N$31881 N$31882 "Straight Waveguide" sch_x=197 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15942 N$31883 N$31884 "Straight Waveguide" sch_x=197 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15943 N$31885 N$31886 "Straight Waveguide" sch_x=197 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15944 N$31887 N$31888 "Straight Waveguide" sch_x=197 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15945 N$31889 N$31890 "Straight Waveguide" sch_x=197 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15946 N$31891 N$31892 "Straight Waveguide" sch_x=197 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15947 N$31893 N$31894 "Straight Waveguide" sch_x=197 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15948 N$31895 N$31896 "Straight Waveguide" sch_x=197 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15949 N$31897 N$31898 "Straight Waveguide" sch_x=197 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15950 N$31899 N$31900 "Straight Waveguide" sch_x=197 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15951 N$31901 N$31902 "Straight Waveguide" sch_x=197 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15952 N$31903 N$31904 "Straight Waveguide" sch_x=197 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15953 N$31905 N$31906 "Straight Waveguide" sch_x=197 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15954 N$31907 N$31908 "Straight Waveguide" sch_x=197 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15955 N$31909 N$31910 "Straight Waveguide" sch_x=197 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15956 N$31911 N$31912 "Straight Waveguide" sch_x=197 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15957 N$31913 N$31914 "Straight Waveguide" sch_x=197 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15958 N$31915 N$31916 "Straight Waveguide" sch_x=197 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15959 N$31917 N$31918 "Straight Waveguide" sch_x=197 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15960 N$31919 N$31920 "Straight Waveguide" sch_x=197 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15961 N$31921 N$31922 "Straight Waveguide" sch_x=197 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15962 N$31923 N$31924 "Straight Waveguide" sch_x=197 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15963 N$31925 N$31926 "Straight Waveguide" sch_x=195 sch_y=33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15964 N$31927 N$31928 "Straight Waveguide" sch_x=195 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15965 N$31929 N$31930 "Straight Waveguide" sch_x=195 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15966 N$31931 N$31932 "Straight Waveguide" sch_x=195 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15967 N$31933 N$31934 "Straight Waveguide" sch_x=195 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15968 N$31935 N$31936 "Straight Waveguide" sch_x=195 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15969 N$31937 N$31938 "Straight Waveguide" sch_x=195 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15970 N$31939 N$31940 "Straight Waveguide" sch_x=195 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15971 N$31941 N$31942 "Straight Waveguide" sch_x=195 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15972 N$31943 N$31944 "Straight Waveguide" sch_x=195 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15973 N$31945 N$31946 "Straight Waveguide" sch_x=195 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15974 N$31947 N$31948 "Straight Waveguide" sch_x=195 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15975 N$31949 N$31950 "Straight Waveguide" sch_x=195 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15976 N$31951 N$31952 "Straight Waveguide" sch_x=195 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15977 N$31953 N$31954 "Straight Waveguide" sch_x=195 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15978 N$31955 N$31956 "Straight Waveguide" sch_x=195 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15979 N$31957 N$31958 "Straight Waveguide" sch_x=195 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15980 N$31959 N$31960 "Straight Waveguide" sch_x=195 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15981 N$31961 N$31962 "Straight Waveguide" sch_x=195 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15982 N$31963 N$31964 "Straight Waveguide" sch_x=195 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15983 N$31965 N$31966 "Straight Waveguide" sch_x=195 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15984 N$31967 N$31968 "Straight Waveguide" sch_x=195 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15985 N$31969 N$31970 "Straight Waveguide" sch_x=195 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15986 N$31971 N$31972 "Straight Waveguide" sch_x=195 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15987 N$31973 N$31974 "Straight Waveguide" sch_x=195 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15988 N$31975 N$31976 "Straight Waveguide" sch_x=195 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15989 N$31977 N$31978 "Straight Waveguide" sch_x=195 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15990 N$31979 N$31980 "Straight Waveguide" sch_x=195 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15991 N$31981 N$31982 "Straight Waveguide" sch_x=195 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15992 N$31983 N$31984 "Straight Waveguide" sch_x=195 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15993 N$31985 N$31986 "Straight Waveguide" sch_x=195 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15994 N$31987 N$31988 "Straight Waveguide" sch_x=195 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15995 N$31989 N$31990 "Straight Waveguide" sch_x=195 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15996 N$31991 N$31992 "Straight Waveguide" sch_x=195 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15997 N$31993 N$31994 "Straight Waveguide" sch_x=195 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15998 N$31995 N$31996 "Straight Waveguide" sch_x=195 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15999 N$31997 N$31998 "Straight Waveguide" sch_x=195 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16000 N$31999 N$32000 "Straight Waveguide" sch_x=195 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16001 N$32001 N$32002 "Straight Waveguide" sch_x=195 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16002 N$32003 N$32004 "Straight Waveguide" sch_x=195 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16003 N$32005 N$32006 "Straight Waveguide" sch_x=195 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16004 N$32007 N$32008 "Straight Waveguide" sch_x=195 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16005 N$32009 N$32010 "Straight Waveguide" sch_x=195 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16006 N$32011 N$32012 "Straight Waveguide" sch_x=195 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16007 N$32013 N$32014 "Straight Waveguide" sch_x=195 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16008 N$32015 N$32016 "Straight Waveguide" sch_x=195 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16009 N$32017 N$32018 "Straight Waveguide" sch_x=195 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16010 N$32019 N$32020 "Straight Waveguide" sch_x=195 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16011 N$32021 N$32022 "Straight Waveguide" sch_x=195 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16012 N$32023 N$32024 "Straight Waveguide" sch_x=195 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16013 N$32025 N$32026 "Straight Waveguide" sch_x=195 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16014 N$32027 N$32028 "Straight Waveguide" sch_x=195 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16015 N$32029 N$32030 "Straight Waveguide" sch_x=195 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16016 N$32031 N$32032 "Straight Waveguide" sch_x=195 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16017 N$32033 N$32034 "Straight Waveguide" sch_x=195 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16018 N$32035 N$32036 "Straight Waveguide" sch_x=195 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16019 N$32037 N$32038 "Straight Waveguide" sch_x=195 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16020 N$32039 N$32040 "Straight Waveguide" sch_x=195 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16021 N$32041 N$32042 "Straight Waveguide" sch_x=195 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16022 N$32043 N$32044 "Straight Waveguide" sch_x=195 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16023 N$32045 N$32046 "Straight Waveguide" sch_x=195 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16024 N$32047 N$32048 "Straight Waveguide" sch_x=195 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16025 N$32049 N$32050 "Straight Waveguide" sch_x=195 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16026 N$32051 N$32052 "Straight Waveguide" sch_x=195 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16027 N$32053 N$32054 "Straight Waveguide" sch_x=195 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16028 N$32055 N$32056 "Straight Waveguide" sch_x=195 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16029 N$32057 N$32058 "Straight Waveguide" sch_x=195 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16030 N$32059 N$32060 "Straight Waveguide" sch_x=195 sch_y=-33.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16031 N$32061 N$32062 "Straight Waveguide" sch_x=193 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16032 N$32063 N$32064 "Straight Waveguide" sch_x=193 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16033 N$32065 N$32066 "Straight Waveguide" sch_x=193 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16034 N$32067 N$32068 "Straight Waveguide" sch_x=193 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16035 N$32069 N$32070 "Straight Waveguide" sch_x=193 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16036 N$32071 N$32072 "Straight Waveguide" sch_x=193 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16037 N$32073 N$32074 "Straight Waveguide" sch_x=193 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16038 N$32075 N$32076 "Straight Waveguide" sch_x=193 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16039 N$32077 N$32078 "Straight Waveguide" sch_x=193 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16040 N$32079 N$32080 "Straight Waveguide" sch_x=193 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16041 N$32081 N$32082 "Straight Waveguide" sch_x=193 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16042 N$32083 N$32084 "Straight Waveguide" sch_x=193 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16043 N$32085 N$32086 "Straight Waveguide" sch_x=193 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16044 N$32087 N$32088 "Straight Waveguide" sch_x=193 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16045 N$32089 N$32090 "Straight Waveguide" sch_x=193 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16046 N$32091 N$32092 "Straight Waveguide" sch_x=193 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16047 N$32093 N$32094 "Straight Waveguide" sch_x=193 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16048 N$32095 N$32096 "Straight Waveguide" sch_x=193 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16049 N$32097 N$32098 "Straight Waveguide" sch_x=193 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16050 N$32099 N$32100 "Straight Waveguide" sch_x=193 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16051 N$32101 N$32102 "Straight Waveguide" sch_x=193 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16052 N$32103 N$32104 "Straight Waveguide" sch_x=193 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16053 N$32105 N$32106 "Straight Waveguide" sch_x=193 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16054 N$32107 N$32108 "Straight Waveguide" sch_x=193 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16055 N$32109 N$32110 "Straight Waveguide" sch_x=193 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16056 N$32111 N$32112 "Straight Waveguide" sch_x=193 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16057 N$32113 N$32114 "Straight Waveguide" sch_x=193 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16058 N$32115 N$32116 "Straight Waveguide" sch_x=193 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16059 N$32117 N$32118 "Straight Waveguide" sch_x=193 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16060 N$32119 N$32120 "Straight Waveguide" sch_x=193 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16061 N$32121 N$32122 "Straight Waveguide" sch_x=193 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16062 N$32123 N$32124 "Straight Waveguide" sch_x=193 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16063 N$32125 N$32126 "Straight Waveguide" sch_x=193 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16064 N$32127 N$32128 "Straight Waveguide" sch_x=193 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16065 N$32129 N$32130 "Straight Waveguide" sch_x=193 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16066 N$32131 N$32132 "Straight Waveguide" sch_x=193 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16067 N$32133 N$32134 "Straight Waveguide" sch_x=193 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16068 N$32135 N$32136 "Straight Waveguide" sch_x=193 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16069 N$32137 N$32138 "Straight Waveguide" sch_x=193 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16070 N$32139 N$32140 "Straight Waveguide" sch_x=193 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16071 N$32141 N$32142 "Straight Waveguide" sch_x=193 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16072 N$32143 N$32144 "Straight Waveguide" sch_x=193 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16073 N$32145 N$32146 "Straight Waveguide" sch_x=193 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16074 N$32147 N$32148 "Straight Waveguide" sch_x=193 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16075 N$32149 N$32150 "Straight Waveguide" sch_x=193 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16076 N$32151 N$32152 "Straight Waveguide" sch_x=193 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16077 N$32153 N$32154 "Straight Waveguide" sch_x=193 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16078 N$32155 N$32156 "Straight Waveguide" sch_x=193 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16079 N$32157 N$32158 "Straight Waveguide" sch_x=193 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16080 N$32159 N$32160 "Straight Waveguide" sch_x=193 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16081 N$32161 N$32162 "Straight Waveguide" sch_x=193 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16082 N$32163 N$32164 "Straight Waveguide" sch_x=193 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16083 N$32165 N$32166 "Straight Waveguide" sch_x=193 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16084 N$32167 N$32168 "Straight Waveguide" sch_x=193 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16085 N$32169 N$32170 "Straight Waveguide" sch_x=193 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16086 N$32171 N$32172 "Straight Waveguide" sch_x=193 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16087 N$32173 N$32174 "Straight Waveguide" sch_x=193 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16088 N$32175 N$32176 "Straight Waveguide" sch_x=193 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16089 N$32177 N$32178 "Straight Waveguide" sch_x=193 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16090 N$32179 N$32180 "Straight Waveguide" sch_x=193 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16091 N$32181 N$32182 "Straight Waveguide" sch_x=193 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16092 N$32183 N$32184 "Straight Waveguide" sch_x=193 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16093 N$32185 N$32186 "Straight Waveguide" sch_x=193 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16094 N$32187 N$32188 "Straight Waveguide" sch_x=193 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16095 N$32189 N$32190 "Straight Waveguide" sch_x=193 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16096 N$32191 N$32192 "Straight Waveguide" sch_x=193 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16097 N$32193 N$32194 "Straight Waveguide" sch_x=191 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16098 N$32195 N$32196 "Straight Waveguide" sch_x=191 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16099 N$32197 N$32198 "Straight Waveguide" sch_x=191 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16100 N$32199 N$32200 "Straight Waveguide" sch_x=191 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16101 N$32201 N$32202 "Straight Waveguide" sch_x=191 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16102 N$32203 N$32204 "Straight Waveguide" sch_x=191 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16103 N$32205 N$32206 "Straight Waveguide" sch_x=191 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16104 N$32207 N$32208 "Straight Waveguide" sch_x=191 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16105 N$32209 N$32210 "Straight Waveguide" sch_x=191 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16106 N$32211 N$32212 "Straight Waveguide" sch_x=191 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16107 N$32213 N$32214 "Straight Waveguide" sch_x=191 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16108 N$32215 N$32216 "Straight Waveguide" sch_x=191 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16109 N$32217 N$32218 "Straight Waveguide" sch_x=191 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16110 N$32219 N$32220 "Straight Waveguide" sch_x=191 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16111 N$32221 N$32222 "Straight Waveguide" sch_x=191 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16112 N$32223 N$32224 "Straight Waveguide" sch_x=191 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16113 N$32225 N$32226 "Straight Waveguide" sch_x=191 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16114 N$32227 N$32228 "Straight Waveguide" sch_x=191 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16115 N$32229 N$32230 "Straight Waveguide" sch_x=191 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16116 N$32231 N$32232 "Straight Waveguide" sch_x=191 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16117 N$32233 N$32234 "Straight Waveguide" sch_x=191 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16118 N$32235 N$32236 "Straight Waveguide" sch_x=191 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16119 N$32237 N$32238 "Straight Waveguide" sch_x=191 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16120 N$32239 N$32240 "Straight Waveguide" sch_x=191 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16121 N$32241 N$32242 "Straight Waveguide" sch_x=191 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16122 N$32243 N$32244 "Straight Waveguide" sch_x=191 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16123 N$32245 N$32246 "Straight Waveguide" sch_x=191 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16124 N$32247 N$32248 "Straight Waveguide" sch_x=191 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16125 N$32249 N$32250 "Straight Waveguide" sch_x=191 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16126 N$32251 N$32252 "Straight Waveguide" sch_x=191 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16127 N$32253 N$32254 "Straight Waveguide" sch_x=191 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16128 N$32255 N$32256 "Straight Waveguide" sch_x=191 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16129 N$32257 N$32258 "Straight Waveguide" sch_x=191 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16130 N$32259 N$32260 "Straight Waveguide" sch_x=191 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16131 N$32261 N$32262 "Straight Waveguide" sch_x=191 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16132 N$32263 N$32264 "Straight Waveguide" sch_x=191 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16133 N$32265 N$32266 "Straight Waveguide" sch_x=191 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16134 N$32267 N$32268 "Straight Waveguide" sch_x=191 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16135 N$32269 N$32270 "Straight Waveguide" sch_x=191 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16136 N$32271 N$32272 "Straight Waveguide" sch_x=191 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16137 N$32273 N$32274 "Straight Waveguide" sch_x=191 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16138 N$32275 N$32276 "Straight Waveguide" sch_x=191 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16139 N$32277 N$32278 "Straight Waveguide" sch_x=191 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16140 N$32279 N$32280 "Straight Waveguide" sch_x=191 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16141 N$32281 N$32282 "Straight Waveguide" sch_x=191 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16142 N$32283 N$32284 "Straight Waveguide" sch_x=191 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16143 N$32285 N$32286 "Straight Waveguide" sch_x=191 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16144 N$32287 N$32288 "Straight Waveguide" sch_x=191 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16145 N$32289 N$32290 "Straight Waveguide" sch_x=191 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16146 N$32291 N$32292 "Straight Waveguide" sch_x=191 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16147 N$32293 N$32294 "Straight Waveguide" sch_x=191 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16148 N$32295 N$32296 "Straight Waveguide" sch_x=191 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16149 N$32297 N$32298 "Straight Waveguide" sch_x=191 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16150 N$32299 N$32300 "Straight Waveguide" sch_x=191 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16151 N$32301 N$32302 "Straight Waveguide" sch_x=191 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16152 N$32303 N$32304 "Straight Waveguide" sch_x=191 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16153 N$32305 N$32306 "Straight Waveguide" sch_x=191 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16154 N$32307 N$32308 "Straight Waveguide" sch_x=191 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16155 N$32309 N$32310 "Straight Waveguide" sch_x=191 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16156 N$32311 N$32312 "Straight Waveguide" sch_x=191 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16157 N$32313 N$32314 "Straight Waveguide" sch_x=191 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16158 N$32315 N$32316 "Straight Waveguide" sch_x=191 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16159 N$32317 N$32318 "Straight Waveguide" sch_x=191 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16160 N$32319 N$32320 "Straight Waveguide" sch_x=191 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16161 N$32321 N$32322 "Straight Waveguide" sch_x=189 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16162 N$32323 N$32324 "Straight Waveguide" sch_x=189 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16163 N$32325 N$32326 "Straight Waveguide" sch_x=189 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16164 N$32327 N$32328 "Straight Waveguide" sch_x=189 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16165 N$32329 N$32330 "Straight Waveguide" sch_x=189 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16166 N$32331 N$32332 "Straight Waveguide" sch_x=189 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16167 N$32333 N$32334 "Straight Waveguide" sch_x=189 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16168 N$32335 N$32336 "Straight Waveguide" sch_x=189 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16169 N$32337 N$32338 "Straight Waveguide" sch_x=189 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16170 N$32339 N$32340 "Straight Waveguide" sch_x=189 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16171 N$32341 N$32342 "Straight Waveguide" sch_x=189 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16172 N$32343 N$32344 "Straight Waveguide" sch_x=189 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16173 N$32345 N$32346 "Straight Waveguide" sch_x=189 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16174 N$32347 N$32348 "Straight Waveguide" sch_x=189 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16175 N$32349 N$32350 "Straight Waveguide" sch_x=189 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16176 N$32351 N$32352 "Straight Waveguide" sch_x=189 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16177 N$32353 N$32354 "Straight Waveguide" sch_x=189 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16178 N$32355 N$32356 "Straight Waveguide" sch_x=189 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16179 N$32357 N$32358 "Straight Waveguide" sch_x=189 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16180 N$32359 N$32360 "Straight Waveguide" sch_x=189 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16181 N$32361 N$32362 "Straight Waveguide" sch_x=189 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16182 N$32363 N$32364 "Straight Waveguide" sch_x=189 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16183 N$32365 N$32366 "Straight Waveguide" sch_x=189 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16184 N$32367 N$32368 "Straight Waveguide" sch_x=189 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16185 N$32369 N$32370 "Straight Waveguide" sch_x=189 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16186 N$32371 N$32372 "Straight Waveguide" sch_x=189 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16187 N$32373 N$32374 "Straight Waveguide" sch_x=189 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16188 N$32375 N$32376 "Straight Waveguide" sch_x=189 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16189 N$32377 N$32378 "Straight Waveguide" sch_x=189 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16190 N$32379 N$32380 "Straight Waveguide" sch_x=189 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16191 N$32381 N$32382 "Straight Waveguide" sch_x=189 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16192 N$32383 N$32384 "Straight Waveguide" sch_x=189 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16193 N$32385 N$32386 "Straight Waveguide" sch_x=189 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16194 N$32387 N$32388 "Straight Waveguide" sch_x=189 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16195 N$32389 N$32390 "Straight Waveguide" sch_x=189 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16196 N$32391 N$32392 "Straight Waveguide" sch_x=189 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16197 N$32393 N$32394 "Straight Waveguide" sch_x=189 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16198 N$32395 N$32396 "Straight Waveguide" sch_x=189 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16199 N$32397 N$32398 "Straight Waveguide" sch_x=189 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16200 N$32399 N$32400 "Straight Waveguide" sch_x=189 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16201 N$32401 N$32402 "Straight Waveguide" sch_x=189 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16202 N$32403 N$32404 "Straight Waveguide" sch_x=189 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16203 N$32405 N$32406 "Straight Waveguide" sch_x=189 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16204 N$32407 N$32408 "Straight Waveguide" sch_x=189 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16205 N$32409 N$32410 "Straight Waveguide" sch_x=189 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16206 N$32411 N$32412 "Straight Waveguide" sch_x=189 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16207 N$32413 N$32414 "Straight Waveguide" sch_x=189 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16208 N$32415 N$32416 "Straight Waveguide" sch_x=189 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16209 N$32417 N$32418 "Straight Waveguide" sch_x=189 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16210 N$32419 N$32420 "Straight Waveguide" sch_x=189 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16211 N$32421 N$32422 "Straight Waveguide" sch_x=189 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16212 N$32423 N$32424 "Straight Waveguide" sch_x=189 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16213 N$32425 N$32426 "Straight Waveguide" sch_x=189 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16214 N$32427 N$32428 "Straight Waveguide" sch_x=189 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16215 N$32429 N$32430 "Straight Waveguide" sch_x=189 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16216 N$32431 N$32432 "Straight Waveguide" sch_x=189 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16217 N$32433 N$32434 "Straight Waveguide" sch_x=189 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16218 N$32435 N$32436 "Straight Waveguide" sch_x=189 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16219 N$32437 N$32438 "Straight Waveguide" sch_x=189 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16220 N$32439 N$32440 "Straight Waveguide" sch_x=189 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16221 N$32441 N$32442 "Straight Waveguide" sch_x=189 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16222 N$32443 N$32444 "Straight Waveguide" sch_x=189 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16223 N$32445 N$32446 "Straight Waveguide" sch_x=187 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16224 N$32447 N$32448 "Straight Waveguide" sch_x=187 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16225 N$32449 N$32450 "Straight Waveguide" sch_x=187 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16226 N$32451 N$32452 "Straight Waveguide" sch_x=187 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16227 N$32453 N$32454 "Straight Waveguide" sch_x=187 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16228 N$32455 N$32456 "Straight Waveguide" sch_x=187 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16229 N$32457 N$32458 "Straight Waveguide" sch_x=187 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16230 N$32459 N$32460 "Straight Waveguide" sch_x=187 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16231 N$32461 N$32462 "Straight Waveguide" sch_x=187 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16232 N$32463 N$32464 "Straight Waveguide" sch_x=187 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16233 N$32465 N$32466 "Straight Waveguide" sch_x=187 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16234 N$32467 N$32468 "Straight Waveguide" sch_x=187 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16235 N$32469 N$32470 "Straight Waveguide" sch_x=187 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16236 N$32471 N$32472 "Straight Waveguide" sch_x=187 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16237 N$32473 N$32474 "Straight Waveguide" sch_x=187 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16238 N$32475 N$32476 "Straight Waveguide" sch_x=187 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16239 N$32477 N$32478 "Straight Waveguide" sch_x=187 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16240 N$32479 N$32480 "Straight Waveguide" sch_x=187 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16241 N$32481 N$32482 "Straight Waveguide" sch_x=187 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16242 N$32483 N$32484 "Straight Waveguide" sch_x=187 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16243 N$32485 N$32486 "Straight Waveguide" sch_x=187 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16244 N$32487 N$32488 "Straight Waveguide" sch_x=187 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16245 N$32489 N$32490 "Straight Waveguide" sch_x=187 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16246 N$32491 N$32492 "Straight Waveguide" sch_x=187 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16247 N$32493 N$32494 "Straight Waveguide" sch_x=187 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16248 N$32495 N$32496 "Straight Waveguide" sch_x=187 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16249 N$32497 N$32498 "Straight Waveguide" sch_x=187 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16250 N$32499 N$32500 "Straight Waveguide" sch_x=187 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16251 N$32501 N$32502 "Straight Waveguide" sch_x=187 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16252 N$32503 N$32504 "Straight Waveguide" sch_x=187 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16253 N$32505 N$32506 "Straight Waveguide" sch_x=187 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16254 N$32507 N$32508 "Straight Waveguide" sch_x=187 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16255 N$32509 N$32510 "Straight Waveguide" sch_x=187 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16256 N$32511 N$32512 "Straight Waveguide" sch_x=187 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16257 N$32513 N$32514 "Straight Waveguide" sch_x=187 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16258 N$32515 N$32516 "Straight Waveguide" sch_x=187 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16259 N$32517 N$32518 "Straight Waveguide" sch_x=187 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16260 N$32519 N$32520 "Straight Waveguide" sch_x=187 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16261 N$32521 N$32522 "Straight Waveguide" sch_x=187 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16262 N$32523 N$32524 "Straight Waveguide" sch_x=187 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16263 N$32525 N$32526 "Straight Waveguide" sch_x=187 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16264 N$32527 N$32528 "Straight Waveguide" sch_x=187 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16265 N$32529 N$32530 "Straight Waveguide" sch_x=187 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16266 N$32531 N$32532 "Straight Waveguide" sch_x=187 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16267 N$32533 N$32534 "Straight Waveguide" sch_x=187 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16268 N$32535 N$32536 "Straight Waveguide" sch_x=187 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16269 N$32537 N$32538 "Straight Waveguide" sch_x=187 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16270 N$32539 N$32540 "Straight Waveguide" sch_x=187 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16271 N$32541 N$32542 "Straight Waveguide" sch_x=187 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16272 N$32543 N$32544 "Straight Waveguide" sch_x=187 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16273 N$32545 N$32546 "Straight Waveguide" sch_x=187 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16274 N$32547 N$32548 "Straight Waveguide" sch_x=187 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16275 N$32549 N$32550 "Straight Waveguide" sch_x=187 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16276 N$32551 N$32552 "Straight Waveguide" sch_x=187 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16277 N$32553 N$32554 "Straight Waveguide" sch_x=187 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16278 N$32555 N$32556 "Straight Waveguide" sch_x=187 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16279 N$32557 N$32558 "Straight Waveguide" sch_x=187 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16280 N$32559 N$32560 "Straight Waveguide" sch_x=187 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16281 N$32561 N$32562 "Straight Waveguide" sch_x=187 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16282 N$32563 N$32564 "Straight Waveguide" sch_x=187 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16283 N$32565 N$32566 "Straight Waveguide" sch_x=185 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16284 N$32567 N$32568 "Straight Waveguide" sch_x=185 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16285 N$32569 N$32570 "Straight Waveguide" sch_x=185 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16286 N$32571 N$32572 "Straight Waveguide" sch_x=185 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16287 N$32573 N$32574 "Straight Waveguide" sch_x=185 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16288 N$32575 N$32576 "Straight Waveguide" sch_x=185 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16289 N$32577 N$32578 "Straight Waveguide" sch_x=185 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16290 N$32579 N$32580 "Straight Waveguide" sch_x=185 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16291 N$32581 N$32582 "Straight Waveguide" sch_x=185 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16292 N$32583 N$32584 "Straight Waveguide" sch_x=185 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16293 N$32585 N$32586 "Straight Waveguide" sch_x=185 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16294 N$32587 N$32588 "Straight Waveguide" sch_x=185 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16295 N$32589 N$32590 "Straight Waveguide" sch_x=185 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16296 N$32591 N$32592 "Straight Waveguide" sch_x=185 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16297 N$32593 N$32594 "Straight Waveguide" sch_x=185 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16298 N$32595 N$32596 "Straight Waveguide" sch_x=185 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16299 N$32597 N$32598 "Straight Waveguide" sch_x=185 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16300 N$32599 N$32600 "Straight Waveguide" sch_x=185 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16301 N$32601 N$32602 "Straight Waveguide" sch_x=185 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16302 N$32603 N$32604 "Straight Waveguide" sch_x=185 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16303 N$32605 N$32606 "Straight Waveguide" sch_x=185 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16304 N$32607 N$32608 "Straight Waveguide" sch_x=185 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16305 N$32609 N$32610 "Straight Waveguide" sch_x=185 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16306 N$32611 N$32612 "Straight Waveguide" sch_x=185 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16307 N$32613 N$32614 "Straight Waveguide" sch_x=185 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16308 N$32615 N$32616 "Straight Waveguide" sch_x=185 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16309 N$32617 N$32618 "Straight Waveguide" sch_x=185 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16310 N$32619 N$32620 "Straight Waveguide" sch_x=185 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16311 N$32621 N$32622 "Straight Waveguide" sch_x=185 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16312 N$32623 N$32624 "Straight Waveguide" sch_x=185 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16313 N$32625 N$32626 "Straight Waveguide" sch_x=185 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16314 N$32627 N$32628 "Straight Waveguide" sch_x=185 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16315 N$32629 N$32630 "Straight Waveguide" sch_x=185 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16316 N$32631 N$32632 "Straight Waveguide" sch_x=185 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16317 N$32633 N$32634 "Straight Waveguide" sch_x=185 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16318 N$32635 N$32636 "Straight Waveguide" sch_x=185 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16319 N$32637 N$32638 "Straight Waveguide" sch_x=185 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16320 N$32639 N$32640 "Straight Waveguide" sch_x=185 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16321 N$32641 N$32642 "Straight Waveguide" sch_x=185 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16322 N$32643 N$32644 "Straight Waveguide" sch_x=185 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16323 N$32645 N$32646 "Straight Waveguide" sch_x=185 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16324 N$32647 N$32648 "Straight Waveguide" sch_x=185 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16325 N$32649 N$32650 "Straight Waveguide" sch_x=185 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16326 N$32651 N$32652 "Straight Waveguide" sch_x=185 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16327 N$32653 N$32654 "Straight Waveguide" sch_x=185 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16328 N$32655 N$32656 "Straight Waveguide" sch_x=185 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16329 N$32657 N$32658 "Straight Waveguide" sch_x=185 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16330 N$32659 N$32660 "Straight Waveguide" sch_x=185 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16331 N$32661 N$32662 "Straight Waveguide" sch_x=185 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16332 N$32663 N$32664 "Straight Waveguide" sch_x=185 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16333 N$32665 N$32666 "Straight Waveguide" sch_x=185 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16334 N$32667 N$32668 "Straight Waveguide" sch_x=185 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16335 N$32669 N$32670 "Straight Waveguide" sch_x=185 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16336 N$32671 N$32672 "Straight Waveguide" sch_x=185 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16337 N$32673 N$32674 "Straight Waveguide" sch_x=185 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16338 N$32675 N$32676 "Straight Waveguide" sch_x=185 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16339 N$32677 N$32678 "Straight Waveguide" sch_x=185 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16340 N$32679 N$32680 "Straight Waveguide" sch_x=185 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16341 N$32681 N$32682 "Straight Waveguide" sch_x=183 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16342 N$32683 N$32684 "Straight Waveguide" sch_x=183 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16343 N$32685 N$32686 "Straight Waveguide" sch_x=183 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16344 N$32687 N$32688 "Straight Waveguide" sch_x=183 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16345 N$32689 N$32690 "Straight Waveguide" sch_x=183 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16346 N$32691 N$32692 "Straight Waveguide" sch_x=183 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16347 N$32693 N$32694 "Straight Waveguide" sch_x=183 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16348 N$32695 N$32696 "Straight Waveguide" sch_x=183 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16349 N$32697 N$32698 "Straight Waveguide" sch_x=183 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16350 N$32699 N$32700 "Straight Waveguide" sch_x=183 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16351 N$32701 N$32702 "Straight Waveguide" sch_x=183 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16352 N$32703 N$32704 "Straight Waveguide" sch_x=183 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16353 N$32705 N$32706 "Straight Waveguide" sch_x=183 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16354 N$32707 N$32708 "Straight Waveguide" sch_x=183 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16355 N$32709 N$32710 "Straight Waveguide" sch_x=183 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16356 N$32711 N$32712 "Straight Waveguide" sch_x=183 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16357 N$32713 N$32714 "Straight Waveguide" sch_x=183 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16358 N$32715 N$32716 "Straight Waveguide" sch_x=183 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16359 N$32717 N$32718 "Straight Waveguide" sch_x=183 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16360 N$32719 N$32720 "Straight Waveguide" sch_x=183 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16361 N$32721 N$32722 "Straight Waveguide" sch_x=183 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16362 N$32723 N$32724 "Straight Waveguide" sch_x=183 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16363 N$32725 N$32726 "Straight Waveguide" sch_x=183 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16364 N$32727 N$32728 "Straight Waveguide" sch_x=183 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16365 N$32729 N$32730 "Straight Waveguide" sch_x=183 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16366 N$32731 N$32732 "Straight Waveguide" sch_x=183 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16367 N$32733 N$32734 "Straight Waveguide" sch_x=183 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16368 N$32735 N$32736 "Straight Waveguide" sch_x=183 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16369 N$32737 N$32738 "Straight Waveguide" sch_x=183 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16370 N$32739 N$32740 "Straight Waveguide" sch_x=183 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16371 N$32741 N$32742 "Straight Waveguide" sch_x=183 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16372 N$32743 N$32744 "Straight Waveguide" sch_x=183 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16373 N$32745 N$32746 "Straight Waveguide" sch_x=183 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16374 N$32747 N$32748 "Straight Waveguide" sch_x=183 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16375 N$32749 N$32750 "Straight Waveguide" sch_x=183 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16376 N$32751 N$32752 "Straight Waveguide" sch_x=183 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16377 N$32753 N$32754 "Straight Waveguide" sch_x=183 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16378 N$32755 N$32756 "Straight Waveguide" sch_x=183 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16379 N$32757 N$32758 "Straight Waveguide" sch_x=183 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16380 N$32759 N$32760 "Straight Waveguide" sch_x=183 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16381 N$32761 N$32762 "Straight Waveguide" sch_x=183 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16382 N$32763 N$32764 "Straight Waveguide" sch_x=183 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16383 N$32765 N$32766 "Straight Waveguide" sch_x=183 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16384 N$32767 N$32768 "Straight Waveguide" sch_x=183 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16385 N$32769 N$32770 "Straight Waveguide" sch_x=183 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16386 N$32771 N$32772 "Straight Waveguide" sch_x=183 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16387 N$32773 N$32774 "Straight Waveguide" sch_x=183 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16388 N$32775 N$32776 "Straight Waveguide" sch_x=183 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16389 N$32777 N$32778 "Straight Waveguide" sch_x=183 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16390 N$32779 N$32780 "Straight Waveguide" sch_x=183 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16391 N$32781 N$32782 "Straight Waveguide" sch_x=183 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16392 N$32783 N$32784 "Straight Waveguide" sch_x=183 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16393 N$32785 N$32786 "Straight Waveguide" sch_x=183 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16394 N$32787 N$32788 "Straight Waveguide" sch_x=183 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16395 N$32789 N$32790 "Straight Waveguide" sch_x=183 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16396 N$32791 N$32792 "Straight Waveguide" sch_x=183 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16397 N$32793 N$32794 "Straight Waveguide" sch_x=181 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16398 N$32795 N$32796 "Straight Waveguide" sch_x=181 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16399 N$32797 N$32798 "Straight Waveguide" sch_x=181 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16400 N$32799 N$32800 "Straight Waveguide" sch_x=181 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16401 N$32801 N$32802 "Straight Waveguide" sch_x=181 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16402 N$32803 N$32804 "Straight Waveguide" sch_x=181 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16403 N$32805 N$32806 "Straight Waveguide" sch_x=181 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16404 N$32807 N$32808 "Straight Waveguide" sch_x=181 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16405 N$32809 N$32810 "Straight Waveguide" sch_x=181 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16406 N$32811 N$32812 "Straight Waveguide" sch_x=181 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16407 N$32813 N$32814 "Straight Waveguide" sch_x=181 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16408 N$32815 N$32816 "Straight Waveguide" sch_x=181 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16409 N$32817 N$32818 "Straight Waveguide" sch_x=181 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16410 N$32819 N$32820 "Straight Waveguide" sch_x=181 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16411 N$32821 N$32822 "Straight Waveguide" sch_x=181 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16412 N$32823 N$32824 "Straight Waveguide" sch_x=181 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16413 N$32825 N$32826 "Straight Waveguide" sch_x=181 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16414 N$32827 N$32828 "Straight Waveguide" sch_x=181 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16415 N$32829 N$32830 "Straight Waveguide" sch_x=181 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16416 N$32831 N$32832 "Straight Waveguide" sch_x=181 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16417 N$32833 N$32834 "Straight Waveguide" sch_x=181 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16418 N$32835 N$32836 "Straight Waveguide" sch_x=181 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16419 N$32837 N$32838 "Straight Waveguide" sch_x=181 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16420 N$32839 N$32840 "Straight Waveguide" sch_x=181 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16421 N$32841 N$32842 "Straight Waveguide" sch_x=181 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16422 N$32843 N$32844 "Straight Waveguide" sch_x=181 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16423 N$32845 N$32846 "Straight Waveguide" sch_x=181 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16424 N$32847 N$32848 "Straight Waveguide" sch_x=181 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16425 N$32849 N$32850 "Straight Waveguide" sch_x=181 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16426 N$32851 N$32852 "Straight Waveguide" sch_x=181 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16427 N$32853 N$32854 "Straight Waveguide" sch_x=181 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16428 N$32855 N$32856 "Straight Waveguide" sch_x=181 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16429 N$32857 N$32858 "Straight Waveguide" sch_x=181 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16430 N$32859 N$32860 "Straight Waveguide" sch_x=181 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16431 N$32861 N$32862 "Straight Waveguide" sch_x=181 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16432 N$32863 N$32864 "Straight Waveguide" sch_x=181 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16433 N$32865 N$32866 "Straight Waveguide" sch_x=181 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16434 N$32867 N$32868 "Straight Waveguide" sch_x=181 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16435 N$32869 N$32870 "Straight Waveguide" sch_x=181 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16436 N$32871 N$32872 "Straight Waveguide" sch_x=181 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16437 N$32873 N$32874 "Straight Waveguide" sch_x=181 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16438 N$32875 N$32876 "Straight Waveguide" sch_x=181 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16439 N$32877 N$32878 "Straight Waveguide" sch_x=181 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16440 N$32879 N$32880 "Straight Waveguide" sch_x=181 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16441 N$32881 N$32882 "Straight Waveguide" sch_x=181 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16442 N$32883 N$32884 "Straight Waveguide" sch_x=181 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16443 N$32885 N$32886 "Straight Waveguide" sch_x=181 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16444 N$32887 N$32888 "Straight Waveguide" sch_x=181 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16445 N$32889 N$32890 "Straight Waveguide" sch_x=181 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16446 N$32891 N$32892 "Straight Waveguide" sch_x=181 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16447 N$32893 N$32894 "Straight Waveguide" sch_x=181 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16448 N$32895 N$32896 "Straight Waveguide" sch_x=181 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16449 N$32897 N$32898 "Straight Waveguide" sch_x=181 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16450 N$32899 N$32900 "Straight Waveguide" sch_x=181 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16451 N$32901 N$32902 "Straight Waveguide" sch_x=179 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16452 N$32903 N$32904 "Straight Waveguide" sch_x=179 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16453 N$32905 N$32906 "Straight Waveguide" sch_x=179 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16454 N$32907 N$32908 "Straight Waveguide" sch_x=179 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16455 N$32909 N$32910 "Straight Waveguide" sch_x=179 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16456 N$32911 N$32912 "Straight Waveguide" sch_x=179 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16457 N$32913 N$32914 "Straight Waveguide" sch_x=179 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16458 N$32915 N$32916 "Straight Waveguide" sch_x=179 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16459 N$32917 N$32918 "Straight Waveguide" sch_x=179 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16460 N$32919 N$32920 "Straight Waveguide" sch_x=179 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16461 N$32921 N$32922 "Straight Waveguide" sch_x=179 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16462 N$32923 N$32924 "Straight Waveguide" sch_x=179 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16463 N$32925 N$32926 "Straight Waveguide" sch_x=179 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16464 N$32927 N$32928 "Straight Waveguide" sch_x=179 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16465 N$32929 N$32930 "Straight Waveguide" sch_x=179 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16466 N$32931 N$32932 "Straight Waveguide" sch_x=179 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16467 N$32933 N$32934 "Straight Waveguide" sch_x=179 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16468 N$32935 N$32936 "Straight Waveguide" sch_x=179 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16469 N$32937 N$32938 "Straight Waveguide" sch_x=179 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16470 N$32939 N$32940 "Straight Waveguide" sch_x=179 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16471 N$32941 N$32942 "Straight Waveguide" sch_x=179 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16472 N$32943 N$32944 "Straight Waveguide" sch_x=179 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16473 N$32945 N$32946 "Straight Waveguide" sch_x=179 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16474 N$32947 N$32948 "Straight Waveguide" sch_x=179 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16475 N$32949 N$32950 "Straight Waveguide" sch_x=179 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16476 N$32951 N$32952 "Straight Waveguide" sch_x=179 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16477 N$32953 N$32954 "Straight Waveguide" sch_x=179 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16478 N$32955 N$32956 "Straight Waveguide" sch_x=179 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16479 N$32957 N$32958 "Straight Waveguide" sch_x=179 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16480 N$32959 N$32960 "Straight Waveguide" sch_x=179 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16481 N$32961 N$32962 "Straight Waveguide" sch_x=179 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16482 N$32963 N$32964 "Straight Waveguide" sch_x=179 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16483 N$32965 N$32966 "Straight Waveguide" sch_x=179 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16484 N$32967 N$32968 "Straight Waveguide" sch_x=179 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16485 N$32969 N$32970 "Straight Waveguide" sch_x=179 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16486 N$32971 N$32972 "Straight Waveguide" sch_x=179 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16487 N$32973 N$32974 "Straight Waveguide" sch_x=179 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16488 N$32975 N$32976 "Straight Waveguide" sch_x=179 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16489 N$32977 N$32978 "Straight Waveguide" sch_x=179 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16490 N$32979 N$32980 "Straight Waveguide" sch_x=179 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16491 N$32981 N$32982 "Straight Waveguide" sch_x=179 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16492 N$32983 N$32984 "Straight Waveguide" sch_x=179 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16493 N$32985 N$32986 "Straight Waveguide" sch_x=179 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16494 N$32987 N$32988 "Straight Waveguide" sch_x=179 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16495 N$32989 N$32990 "Straight Waveguide" sch_x=179 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16496 N$32991 N$32992 "Straight Waveguide" sch_x=179 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16497 N$32993 N$32994 "Straight Waveguide" sch_x=179 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16498 N$32995 N$32996 "Straight Waveguide" sch_x=179 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16499 N$32997 N$32998 "Straight Waveguide" sch_x=179 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16500 N$32999 N$33000 "Straight Waveguide" sch_x=179 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16501 N$33001 N$33002 "Straight Waveguide" sch_x=179 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16502 N$33003 N$33004 "Straight Waveguide" sch_x=179 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16503 N$33005 N$33006 "Straight Waveguide" sch_x=177 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16504 N$33007 N$33008 "Straight Waveguide" sch_x=177 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16505 N$33009 N$33010 "Straight Waveguide" sch_x=177 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16506 N$33011 N$33012 "Straight Waveguide" sch_x=177 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16507 N$33013 N$33014 "Straight Waveguide" sch_x=177 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16508 N$33015 N$33016 "Straight Waveguide" sch_x=177 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16509 N$33017 N$33018 "Straight Waveguide" sch_x=177 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16510 N$33019 N$33020 "Straight Waveguide" sch_x=177 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16511 N$33021 N$33022 "Straight Waveguide" sch_x=177 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16512 N$33023 N$33024 "Straight Waveguide" sch_x=177 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16513 N$33025 N$33026 "Straight Waveguide" sch_x=177 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16514 N$33027 N$33028 "Straight Waveguide" sch_x=177 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16515 N$33029 N$33030 "Straight Waveguide" sch_x=177 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16516 N$33031 N$33032 "Straight Waveguide" sch_x=177 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16517 N$33033 N$33034 "Straight Waveguide" sch_x=177 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16518 N$33035 N$33036 "Straight Waveguide" sch_x=177 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16519 N$33037 N$33038 "Straight Waveguide" sch_x=177 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16520 N$33039 N$33040 "Straight Waveguide" sch_x=177 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16521 N$33041 N$33042 "Straight Waveguide" sch_x=177 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16522 N$33043 N$33044 "Straight Waveguide" sch_x=177 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16523 N$33045 N$33046 "Straight Waveguide" sch_x=177 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16524 N$33047 N$33048 "Straight Waveguide" sch_x=177 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16525 N$33049 N$33050 "Straight Waveguide" sch_x=177 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16526 N$33051 N$33052 "Straight Waveguide" sch_x=177 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16527 N$33053 N$33054 "Straight Waveguide" sch_x=177 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16528 N$33055 N$33056 "Straight Waveguide" sch_x=177 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16529 N$33057 N$33058 "Straight Waveguide" sch_x=177 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16530 N$33059 N$33060 "Straight Waveguide" sch_x=177 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16531 N$33061 N$33062 "Straight Waveguide" sch_x=177 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16532 N$33063 N$33064 "Straight Waveguide" sch_x=177 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16533 N$33065 N$33066 "Straight Waveguide" sch_x=177 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16534 N$33067 N$33068 "Straight Waveguide" sch_x=177 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16535 N$33069 N$33070 "Straight Waveguide" sch_x=177 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16536 N$33071 N$33072 "Straight Waveguide" sch_x=177 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16537 N$33073 N$33074 "Straight Waveguide" sch_x=177 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16538 N$33075 N$33076 "Straight Waveguide" sch_x=177 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16539 N$33077 N$33078 "Straight Waveguide" sch_x=177 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16540 N$33079 N$33080 "Straight Waveguide" sch_x=177 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16541 N$33081 N$33082 "Straight Waveguide" sch_x=177 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16542 N$33083 N$33084 "Straight Waveguide" sch_x=177 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16543 N$33085 N$33086 "Straight Waveguide" sch_x=177 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16544 N$33087 N$33088 "Straight Waveguide" sch_x=177 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16545 N$33089 N$33090 "Straight Waveguide" sch_x=177 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16546 N$33091 N$33092 "Straight Waveguide" sch_x=177 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16547 N$33093 N$33094 "Straight Waveguide" sch_x=177 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16548 N$33095 N$33096 "Straight Waveguide" sch_x=177 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16549 N$33097 N$33098 "Straight Waveguide" sch_x=177 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16550 N$33099 N$33100 "Straight Waveguide" sch_x=177 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16551 N$33101 N$33102 "Straight Waveguide" sch_x=177 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16552 N$33103 N$33104 "Straight Waveguide" sch_x=177 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16553 N$33105 N$33106 "Straight Waveguide" sch_x=175 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16554 N$33107 N$33108 "Straight Waveguide" sch_x=175 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16555 N$33109 N$33110 "Straight Waveguide" sch_x=175 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16556 N$33111 N$33112 "Straight Waveguide" sch_x=175 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16557 N$33113 N$33114 "Straight Waveguide" sch_x=175 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16558 N$33115 N$33116 "Straight Waveguide" sch_x=175 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16559 N$33117 N$33118 "Straight Waveguide" sch_x=175 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16560 N$33119 N$33120 "Straight Waveguide" sch_x=175 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16561 N$33121 N$33122 "Straight Waveguide" sch_x=175 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16562 N$33123 N$33124 "Straight Waveguide" sch_x=175 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16563 N$33125 N$33126 "Straight Waveguide" sch_x=175 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16564 N$33127 N$33128 "Straight Waveguide" sch_x=175 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16565 N$33129 N$33130 "Straight Waveguide" sch_x=175 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16566 N$33131 N$33132 "Straight Waveguide" sch_x=175 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16567 N$33133 N$33134 "Straight Waveguide" sch_x=175 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16568 N$33135 N$33136 "Straight Waveguide" sch_x=175 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16569 N$33137 N$33138 "Straight Waveguide" sch_x=175 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16570 N$33139 N$33140 "Straight Waveguide" sch_x=175 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16571 N$33141 N$33142 "Straight Waveguide" sch_x=175 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16572 N$33143 N$33144 "Straight Waveguide" sch_x=175 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16573 N$33145 N$33146 "Straight Waveguide" sch_x=175 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16574 N$33147 N$33148 "Straight Waveguide" sch_x=175 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16575 N$33149 N$33150 "Straight Waveguide" sch_x=175 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16576 N$33151 N$33152 "Straight Waveguide" sch_x=175 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16577 N$33153 N$33154 "Straight Waveguide" sch_x=175 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16578 N$33155 N$33156 "Straight Waveguide" sch_x=175 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16579 N$33157 N$33158 "Straight Waveguide" sch_x=175 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16580 N$33159 N$33160 "Straight Waveguide" sch_x=175 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16581 N$33161 N$33162 "Straight Waveguide" sch_x=175 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16582 N$33163 N$33164 "Straight Waveguide" sch_x=175 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16583 N$33165 N$33166 "Straight Waveguide" sch_x=175 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16584 N$33167 N$33168 "Straight Waveguide" sch_x=175 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16585 N$33169 N$33170 "Straight Waveguide" sch_x=175 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16586 N$33171 N$33172 "Straight Waveguide" sch_x=175 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16587 N$33173 N$33174 "Straight Waveguide" sch_x=175 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16588 N$33175 N$33176 "Straight Waveguide" sch_x=175 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16589 N$33177 N$33178 "Straight Waveguide" sch_x=175 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16590 N$33179 N$33180 "Straight Waveguide" sch_x=175 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16591 N$33181 N$33182 "Straight Waveguide" sch_x=175 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16592 N$33183 N$33184 "Straight Waveguide" sch_x=175 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16593 N$33185 N$33186 "Straight Waveguide" sch_x=175 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16594 N$33187 N$33188 "Straight Waveguide" sch_x=175 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16595 N$33189 N$33190 "Straight Waveguide" sch_x=175 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16596 N$33191 N$33192 "Straight Waveguide" sch_x=175 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16597 N$33193 N$33194 "Straight Waveguide" sch_x=175 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16598 N$33195 N$33196 "Straight Waveguide" sch_x=175 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16599 N$33197 N$33198 "Straight Waveguide" sch_x=175 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16600 N$33199 N$33200 "Straight Waveguide" sch_x=175 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16601 N$33201 N$33202 "Straight Waveguide" sch_x=173 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16602 N$33203 N$33204 "Straight Waveguide" sch_x=173 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16603 N$33205 N$33206 "Straight Waveguide" sch_x=173 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16604 N$33207 N$33208 "Straight Waveguide" sch_x=173 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16605 N$33209 N$33210 "Straight Waveguide" sch_x=173 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16606 N$33211 N$33212 "Straight Waveguide" sch_x=173 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16607 N$33213 N$33214 "Straight Waveguide" sch_x=173 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16608 N$33215 N$33216 "Straight Waveguide" sch_x=173 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16609 N$33217 N$33218 "Straight Waveguide" sch_x=173 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16610 N$33219 N$33220 "Straight Waveguide" sch_x=173 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16611 N$33221 N$33222 "Straight Waveguide" sch_x=173 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16612 N$33223 N$33224 "Straight Waveguide" sch_x=173 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16613 N$33225 N$33226 "Straight Waveguide" sch_x=173 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16614 N$33227 N$33228 "Straight Waveguide" sch_x=173 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16615 N$33229 N$33230 "Straight Waveguide" sch_x=173 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16616 N$33231 N$33232 "Straight Waveguide" sch_x=173 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16617 N$33233 N$33234 "Straight Waveguide" sch_x=173 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16618 N$33235 N$33236 "Straight Waveguide" sch_x=173 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16619 N$33237 N$33238 "Straight Waveguide" sch_x=173 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16620 N$33239 N$33240 "Straight Waveguide" sch_x=173 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16621 N$33241 N$33242 "Straight Waveguide" sch_x=173 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16622 N$33243 N$33244 "Straight Waveguide" sch_x=173 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16623 N$33245 N$33246 "Straight Waveguide" sch_x=173 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16624 N$33247 N$33248 "Straight Waveguide" sch_x=173 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16625 N$33249 N$33250 "Straight Waveguide" sch_x=173 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16626 N$33251 N$33252 "Straight Waveguide" sch_x=173 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16627 N$33253 N$33254 "Straight Waveguide" sch_x=173 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16628 N$33255 N$33256 "Straight Waveguide" sch_x=173 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16629 N$33257 N$33258 "Straight Waveguide" sch_x=173 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16630 N$33259 N$33260 "Straight Waveguide" sch_x=173 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16631 N$33261 N$33262 "Straight Waveguide" sch_x=173 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16632 N$33263 N$33264 "Straight Waveguide" sch_x=173 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16633 N$33265 N$33266 "Straight Waveguide" sch_x=173 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16634 N$33267 N$33268 "Straight Waveguide" sch_x=173 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16635 N$33269 N$33270 "Straight Waveguide" sch_x=173 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16636 N$33271 N$33272 "Straight Waveguide" sch_x=173 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16637 N$33273 N$33274 "Straight Waveguide" sch_x=173 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16638 N$33275 N$33276 "Straight Waveguide" sch_x=173 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16639 N$33277 N$33278 "Straight Waveguide" sch_x=173 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16640 N$33279 N$33280 "Straight Waveguide" sch_x=173 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16641 N$33281 N$33282 "Straight Waveguide" sch_x=173 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16642 N$33283 N$33284 "Straight Waveguide" sch_x=173 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16643 N$33285 N$33286 "Straight Waveguide" sch_x=173 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16644 N$33287 N$33288 "Straight Waveguide" sch_x=173 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16645 N$33289 N$33290 "Straight Waveguide" sch_x=173 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16646 N$33291 N$33292 "Straight Waveguide" sch_x=173 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16647 N$33293 N$33294 "Straight Waveguide" sch_x=171 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16648 N$33295 N$33296 "Straight Waveguide" sch_x=171 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16649 N$33297 N$33298 "Straight Waveguide" sch_x=171 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16650 N$33299 N$33300 "Straight Waveguide" sch_x=171 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16651 N$33301 N$33302 "Straight Waveguide" sch_x=171 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16652 N$33303 N$33304 "Straight Waveguide" sch_x=171 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16653 N$33305 N$33306 "Straight Waveguide" sch_x=171 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16654 N$33307 N$33308 "Straight Waveguide" sch_x=171 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16655 N$33309 N$33310 "Straight Waveguide" sch_x=171 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16656 N$33311 N$33312 "Straight Waveguide" sch_x=171 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16657 N$33313 N$33314 "Straight Waveguide" sch_x=171 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16658 N$33315 N$33316 "Straight Waveguide" sch_x=171 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16659 N$33317 N$33318 "Straight Waveguide" sch_x=171 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16660 N$33319 N$33320 "Straight Waveguide" sch_x=171 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16661 N$33321 N$33322 "Straight Waveguide" sch_x=171 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16662 N$33323 N$33324 "Straight Waveguide" sch_x=171 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16663 N$33325 N$33326 "Straight Waveguide" sch_x=171 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16664 N$33327 N$33328 "Straight Waveguide" sch_x=171 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16665 N$33329 N$33330 "Straight Waveguide" sch_x=171 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16666 N$33331 N$33332 "Straight Waveguide" sch_x=171 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16667 N$33333 N$33334 "Straight Waveguide" sch_x=171 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16668 N$33335 N$33336 "Straight Waveguide" sch_x=171 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16669 N$33337 N$33338 "Straight Waveguide" sch_x=171 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16670 N$33339 N$33340 "Straight Waveguide" sch_x=171 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16671 N$33341 N$33342 "Straight Waveguide" sch_x=171 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16672 N$33343 N$33344 "Straight Waveguide" sch_x=171 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16673 N$33345 N$33346 "Straight Waveguide" sch_x=171 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16674 N$33347 N$33348 "Straight Waveguide" sch_x=171 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16675 N$33349 N$33350 "Straight Waveguide" sch_x=171 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16676 N$33351 N$33352 "Straight Waveguide" sch_x=171 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16677 N$33353 N$33354 "Straight Waveguide" sch_x=171 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16678 N$33355 N$33356 "Straight Waveguide" sch_x=171 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16679 N$33357 N$33358 "Straight Waveguide" sch_x=171 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16680 N$33359 N$33360 "Straight Waveguide" sch_x=171 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16681 N$33361 N$33362 "Straight Waveguide" sch_x=171 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16682 N$33363 N$33364 "Straight Waveguide" sch_x=171 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16683 N$33365 N$33366 "Straight Waveguide" sch_x=171 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16684 N$33367 N$33368 "Straight Waveguide" sch_x=171 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16685 N$33369 N$33370 "Straight Waveguide" sch_x=171 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16686 N$33371 N$33372 "Straight Waveguide" sch_x=171 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16687 N$33373 N$33374 "Straight Waveguide" sch_x=171 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16688 N$33375 N$33376 "Straight Waveguide" sch_x=171 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16689 N$33377 N$33378 "Straight Waveguide" sch_x=171 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16690 N$33379 N$33380 "Straight Waveguide" sch_x=171 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16691 N$33381 N$33382 "Straight Waveguide" sch_x=169 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16692 N$33383 N$33384 "Straight Waveguide" sch_x=169 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16693 N$33385 N$33386 "Straight Waveguide" sch_x=169 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16694 N$33387 N$33388 "Straight Waveguide" sch_x=169 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16695 N$33389 N$33390 "Straight Waveguide" sch_x=169 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16696 N$33391 N$33392 "Straight Waveguide" sch_x=169 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16697 N$33393 N$33394 "Straight Waveguide" sch_x=169 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16698 N$33395 N$33396 "Straight Waveguide" sch_x=169 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16699 N$33397 N$33398 "Straight Waveguide" sch_x=169 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16700 N$33399 N$33400 "Straight Waveguide" sch_x=169 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16701 N$33401 N$33402 "Straight Waveguide" sch_x=169 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16702 N$33403 N$33404 "Straight Waveguide" sch_x=169 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16703 N$33405 N$33406 "Straight Waveguide" sch_x=169 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16704 N$33407 N$33408 "Straight Waveguide" sch_x=169 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16705 N$33409 N$33410 "Straight Waveguide" sch_x=169 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16706 N$33411 N$33412 "Straight Waveguide" sch_x=169 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16707 N$33413 N$33414 "Straight Waveguide" sch_x=169 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16708 N$33415 N$33416 "Straight Waveguide" sch_x=169 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16709 N$33417 N$33418 "Straight Waveguide" sch_x=169 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16710 N$33419 N$33420 "Straight Waveguide" sch_x=169 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16711 N$33421 N$33422 "Straight Waveguide" sch_x=169 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16712 N$33423 N$33424 "Straight Waveguide" sch_x=169 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16713 N$33425 N$33426 "Straight Waveguide" sch_x=169 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16714 N$33427 N$33428 "Straight Waveguide" sch_x=169 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16715 N$33429 N$33430 "Straight Waveguide" sch_x=169 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16716 N$33431 N$33432 "Straight Waveguide" sch_x=169 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16717 N$33433 N$33434 "Straight Waveguide" sch_x=169 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16718 N$33435 N$33436 "Straight Waveguide" sch_x=169 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16719 N$33437 N$33438 "Straight Waveguide" sch_x=169 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16720 N$33439 N$33440 "Straight Waveguide" sch_x=169 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16721 N$33441 N$33442 "Straight Waveguide" sch_x=169 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16722 N$33443 N$33444 "Straight Waveguide" sch_x=169 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16723 N$33445 N$33446 "Straight Waveguide" sch_x=169 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16724 N$33447 N$33448 "Straight Waveguide" sch_x=169 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16725 N$33449 N$33450 "Straight Waveguide" sch_x=169 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16726 N$33451 N$33452 "Straight Waveguide" sch_x=169 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16727 N$33453 N$33454 "Straight Waveguide" sch_x=169 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16728 N$33455 N$33456 "Straight Waveguide" sch_x=169 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16729 N$33457 N$33458 "Straight Waveguide" sch_x=169 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16730 N$33459 N$33460 "Straight Waveguide" sch_x=169 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16731 N$33461 N$33462 "Straight Waveguide" sch_x=169 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16732 N$33463 N$33464 "Straight Waveguide" sch_x=169 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16733 N$33465 N$33466 "Straight Waveguide" sch_x=167 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16734 N$33467 N$33468 "Straight Waveguide" sch_x=167 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16735 N$33469 N$33470 "Straight Waveguide" sch_x=167 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16736 N$33471 N$33472 "Straight Waveguide" sch_x=167 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16737 N$33473 N$33474 "Straight Waveguide" sch_x=167 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16738 N$33475 N$33476 "Straight Waveguide" sch_x=167 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16739 N$33477 N$33478 "Straight Waveguide" sch_x=167 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16740 N$33479 N$33480 "Straight Waveguide" sch_x=167 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16741 N$33481 N$33482 "Straight Waveguide" sch_x=167 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16742 N$33483 N$33484 "Straight Waveguide" sch_x=167 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16743 N$33485 N$33486 "Straight Waveguide" sch_x=167 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16744 N$33487 N$33488 "Straight Waveguide" sch_x=167 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16745 N$33489 N$33490 "Straight Waveguide" sch_x=167 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16746 N$33491 N$33492 "Straight Waveguide" sch_x=167 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16747 N$33493 N$33494 "Straight Waveguide" sch_x=167 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16748 N$33495 N$33496 "Straight Waveguide" sch_x=167 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16749 N$33497 N$33498 "Straight Waveguide" sch_x=167 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16750 N$33499 N$33500 "Straight Waveguide" sch_x=167 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16751 N$33501 N$33502 "Straight Waveguide" sch_x=167 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16752 N$33503 N$33504 "Straight Waveguide" sch_x=167 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16753 N$33505 N$33506 "Straight Waveguide" sch_x=167 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16754 N$33507 N$33508 "Straight Waveguide" sch_x=167 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16755 N$33509 N$33510 "Straight Waveguide" sch_x=167 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16756 N$33511 N$33512 "Straight Waveguide" sch_x=167 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16757 N$33513 N$33514 "Straight Waveguide" sch_x=167 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16758 N$33515 N$33516 "Straight Waveguide" sch_x=167 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16759 N$33517 N$33518 "Straight Waveguide" sch_x=167 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16760 N$33519 N$33520 "Straight Waveguide" sch_x=167 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16761 N$33521 N$33522 "Straight Waveguide" sch_x=167 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16762 N$33523 N$33524 "Straight Waveguide" sch_x=167 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16763 N$33525 N$33526 "Straight Waveguide" sch_x=167 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16764 N$33527 N$33528 "Straight Waveguide" sch_x=167 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16765 N$33529 N$33530 "Straight Waveguide" sch_x=167 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16766 N$33531 N$33532 "Straight Waveguide" sch_x=167 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16767 N$33533 N$33534 "Straight Waveguide" sch_x=167 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16768 N$33535 N$33536 "Straight Waveguide" sch_x=167 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16769 N$33537 N$33538 "Straight Waveguide" sch_x=167 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16770 N$33539 N$33540 "Straight Waveguide" sch_x=167 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16771 N$33541 N$33542 "Straight Waveguide" sch_x=167 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16772 N$33543 N$33544 "Straight Waveguide" sch_x=167 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16773 N$33545 N$33546 "Straight Waveguide" sch_x=165 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16774 N$33547 N$33548 "Straight Waveguide" sch_x=165 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16775 N$33549 N$33550 "Straight Waveguide" sch_x=165 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16776 N$33551 N$33552 "Straight Waveguide" sch_x=165 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16777 N$33553 N$33554 "Straight Waveguide" sch_x=165 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16778 N$33555 N$33556 "Straight Waveguide" sch_x=165 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16779 N$33557 N$33558 "Straight Waveguide" sch_x=165 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16780 N$33559 N$33560 "Straight Waveguide" sch_x=165 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16781 N$33561 N$33562 "Straight Waveguide" sch_x=165 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16782 N$33563 N$33564 "Straight Waveguide" sch_x=165 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16783 N$33565 N$33566 "Straight Waveguide" sch_x=165 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16784 N$33567 N$33568 "Straight Waveguide" sch_x=165 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16785 N$33569 N$33570 "Straight Waveguide" sch_x=165 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16786 N$33571 N$33572 "Straight Waveguide" sch_x=165 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16787 N$33573 N$33574 "Straight Waveguide" sch_x=165 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16788 N$33575 N$33576 "Straight Waveguide" sch_x=165 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16789 N$33577 N$33578 "Straight Waveguide" sch_x=165 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16790 N$33579 N$33580 "Straight Waveguide" sch_x=165 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16791 N$33581 N$33582 "Straight Waveguide" sch_x=165 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16792 N$33583 N$33584 "Straight Waveguide" sch_x=165 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16793 N$33585 N$33586 "Straight Waveguide" sch_x=165 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16794 N$33587 N$33588 "Straight Waveguide" sch_x=165 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16795 N$33589 N$33590 "Straight Waveguide" sch_x=165 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16796 N$33591 N$33592 "Straight Waveguide" sch_x=165 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16797 N$33593 N$33594 "Straight Waveguide" sch_x=165 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16798 N$33595 N$33596 "Straight Waveguide" sch_x=165 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16799 N$33597 N$33598 "Straight Waveguide" sch_x=165 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16800 N$33599 N$33600 "Straight Waveguide" sch_x=165 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16801 N$33601 N$33602 "Straight Waveguide" sch_x=165 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16802 N$33603 N$33604 "Straight Waveguide" sch_x=165 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16803 N$33605 N$33606 "Straight Waveguide" sch_x=165 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16804 N$33607 N$33608 "Straight Waveguide" sch_x=165 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16805 N$33609 N$33610 "Straight Waveguide" sch_x=165 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16806 N$33611 N$33612 "Straight Waveguide" sch_x=165 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16807 N$33613 N$33614 "Straight Waveguide" sch_x=165 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16808 N$33615 N$33616 "Straight Waveguide" sch_x=165 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16809 N$33617 N$33618 "Straight Waveguide" sch_x=165 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16810 N$33619 N$33620 "Straight Waveguide" sch_x=165 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16811 N$33621 N$33622 "Straight Waveguide" sch_x=163 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16812 N$33623 N$33624 "Straight Waveguide" sch_x=163 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16813 N$33625 N$33626 "Straight Waveguide" sch_x=163 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16814 N$33627 N$33628 "Straight Waveguide" sch_x=163 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16815 N$33629 N$33630 "Straight Waveguide" sch_x=163 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16816 N$33631 N$33632 "Straight Waveguide" sch_x=163 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16817 N$33633 N$33634 "Straight Waveguide" sch_x=163 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16818 N$33635 N$33636 "Straight Waveguide" sch_x=163 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16819 N$33637 N$33638 "Straight Waveguide" sch_x=163 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16820 N$33639 N$33640 "Straight Waveguide" sch_x=163 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16821 N$33641 N$33642 "Straight Waveguide" sch_x=163 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16822 N$33643 N$33644 "Straight Waveguide" sch_x=163 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16823 N$33645 N$33646 "Straight Waveguide" sch_x=163 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16824 N$33647 N$33648 "Straight Waveguide" sch_x=163 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16825 N$33649 N$33650 "Straight Waveguide" sch_x=163 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16826 N$33651 N$33652 "Straight Waveguide" sch_x=163 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16827 N$33653 N$33654 "Straight Waveguide" sch_x=163 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16828 N$33655 N$33656 "Straight Waveguide" sch_x=163 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16829 N$33657 N$33658 "Straight Waveguide" sch_x=163 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16830 N$33659 N$33660 "Straight Waveguide" sch_x=163 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16831 N$33661 N$33662 "Straight Waveguide" sch_x=163 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16832 N$33663 N$33664 "Straight Waveguide" sch_x=163 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16833 N$33665 N$33666 "Straight Waveguide" sch_x=163 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16834 N$33667 N$33668 "Straight Waveguide" sch_x=163 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16835 N$33669 N$33670 "Straight Waveguide" sch_x=163 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16836 N$33671 N$33672 "Straight Waveguide" sch_x=163 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16837 N$33673 N$33674 "Straight Waveguide" sch_x=163 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16838 N$33675 N$33676 "Straight Waveguide" sch_x=163 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16839 N$33677 N$33678 "Straight Waveguide" sch_x=163 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16840 N$33679 N$33680 "Straight Waveguide" sch_x=163 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16841 N$33681 N$33682 "Straight Waveguide" sch_x=163 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16842 N$33683 N$33684 "Straight Waveguide" sch_x=163 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16843 N$33685 N$33686 "Straight Waveguide" sch_x=163 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16844 N$33687 N$33688 "Straight Waveguide" sch_x=163 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16845 N$33689 N$33690 "Straight Waveguide" sch_x=163 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16846 N$33691 N$33692 "Straight Waveguide" sch_x=163 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16847 N$33693 N$33694 "Straight Waveguide" sch_x=161 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16848 N$33695 N$33696 "Straight Waveguide" sch_x=161 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16849 N$33697 N$33698 "Straight Waveguide" sch_x=161 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16850 N$33699 N$33700 "Straight Waveguide" sch_x=161 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16851 N$33701 N$33702 "Straight Waveguide" sch_x=161 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16852 N$33703 N$33704 "Straight Waveguide" sch_x=161 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16853 N$33705 N$33706 "Straight Waveguide" sch_x=161 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16854 N$33707 N$33708 "Straight Waveguide" sch_x=161 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16855 N$33709 N$33710 "Straight Waveguide" sch_x=161 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16856 N$33711 N$33712 "Straight Waveguide" sch_x=161 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16857 N$33713 N$33714 "Straight Waveguide" sch_x=161 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16858 N$33715 N$33716 "Straight Waveguide" sch_x=161 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16859 N$33717 N$33718 "Straight Waveguide" sch_x=161 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16860 N$33719 N$33720 "Straight Waveguide" sch_x=161 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16861 N$33721 N$33722 "Straight Waveguide" sch_x=161 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16862 N$33723 N$33724 "Straight Waveguide" sch_x=161 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16863 N$33725 N$33726 "Straight Waveguide" sch_x=161 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16864 N$33727 N$33728 "Straight Waveguide" sch_x=161 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16865 N$33729 N$33730 "Straight Waveguide" sch_x=161 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16866 N$33731 N$33732 "Straight Waveguide" sch_x=161 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16867 N$33733 N$33734 "Straight Waveguide" sch_x=161 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16868 N$33735 N$33736 "Straight Waveguide" sch_x=161 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16869 N$33737 N$33738 "Straight Waveguide" sch_x=161 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16870 N$33739 N$33740 "Straight Waveguide" sch_x=161 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16871 N$33741 N$33742 "Straight Waveguide" sch_x=161 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16872 N$33743 N$33744 "Straight Waveguide" sch_x=161 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16873 N$33745 N$33746 "Straight Waveguide" sch_x=161 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16874 N$33747 N$33748 "Straight Waveguide" sch_x=161 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16875 N$33749 N$33750 "Straight Waveguide" sch_x=161 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16876 N$33751 N$33752 "Straight Waveguide" sch_x=161 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16877 N$33753 N$33754 "Straight Waveguide" sch_x=161 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16878 N$33755 N$33756 "Straight Waveguide" sch_x=161 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16879 N$33757 N$33758 "Straight Waveguide" sch_x=161 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16880 N$33759 N$33760 "Straight Waveguide" sch_x=161 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16881 N$33761 N$33762 "Straight Waveguide" sch_x=159 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16882 N$33763 N$33764 "Straight Waveguide" sch_x=159 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16883 N$33765 N$33766 "Straight Waveguide" sch_x=159 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16884 N$33767 N$33768 "Straight Waveguide" sch_x=159 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16885 N$33769 N$33770 "Straight Waveguide" sch_x=159 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16886 N$33771 N$33772 "Straight Waveguide" sch_x=159 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16887 N$33773 N$33774 "Straight Waveguide" sch_x=159 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16888 N$33775 N$33776 "Straight Waveguide" sch_x=159 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16889 N$33777 N$33778 "Straight Waveguide" sch_x=159 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16890 N$33779 N$33780 "Straight Waveguide" sch_x=159 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16891 N$33781 N$33782 "Straight Waveguide" sch_x=159 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16892 N$33783 N$33784 "Straight Waveguide" sch_x=159 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16893 N$33785 N$33786 "Straight Waveguide" sch_x=159 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16894 N$33787 N$33788 "Straight Waveguide" sch_x=159 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16895 N$33789 N$33790 "Straight Waveguide" sch_x=159 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16896 N$33791 N$33792 "Straight Waveguide" sch_x=159 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16897 N$33793 N$33794 "Straight Waveguide" sch_x=159 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16898 N$33795 N$33796 "Straight Waveguide" sch_x=159 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16899 N$33797 N$33798 "Straight Waveguide" sch_x=159 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16900 N$33799 N$33800 "Straight Waveguide" sch_x=159 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16901 N$33801 N$33802 "Straight Waveguide" sch_x=159 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16902 N$33803 N$33804 "Straight Waveguide" sch_x=159 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16903 N$33805 N$33806 "Straight Waveguide" sch_x=159 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16904 N$33807 N$33808 "Straight Waveguide" sch_x=159 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16905 N$33809 N$33810 "Straight Waveguide" sch_x=159 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16906 N$33811 N$33812 "Straight Waveguide" sch_x=159 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16907 N$33813 N$33814 "Straight Waveguide" sch_x=159 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16908 N$33815 N$33816 "Straight Waveguide" sch_x=159 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16909 N$33817 N$33818 "Straight Waveguide" sch_x=159 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16910 N$33819 N$33820 "Straight Waveguide" sch_x=159 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16911 N$33821 N$33822 "Straight Waveguide" sch_x=159 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16912 N$33823 N$33824 "Straight Waveguide" sch_x=159 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16913 N$33825 N$33826 "Straight Waveguide" sch_x=157 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16914 N$33827 N$33828 "Straight Waveguide" sch_x=157 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16915 N$33829 N$33830 "Straight Waveguide" sch_x=157 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16916 N$33831 N$33832 "Straight Waveguide" sch_x=157 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16917 N$33833 N$33834 "Straight Waveguide" sch_x=157 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16918 N$33835 N$33836 "Straight Waveguide" sch_x=157 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16919 N$33837 N$33838 "Straight Waveguide" sch_x=157 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16920 N$33839 N$33840 "Straight Waveguide" sch_x=157 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16921 N$33841 N$33842 "Straight Waveguide" sch_x=157 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16922 N$33843 N$33844 "Straight Waveguide" sch_x=157 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16923 N$33845 N$33846 "Straight Waveguide" sch_x=157 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16924 N$33847 N$33848 "Straight Waveguide" sch_x=157 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16925 N$33849 N$33850 "Straight Waveguide" sch_x=157 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16926 N$33851 N$33852 "Straight Waveguide" sch_x=157 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16927 N$33853 N$33854 "Straight Waveguide" sch_x=157 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16928 N$33855 N$33856 "Straight Waveguide" sch_x=157 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16929 N$33857 N$33858 "Straight Waveguide" sch_x=157 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16930 N$33859 N$33860 "Straight Waveguide" sch_x=157 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16931 N$33861 N$33862 "Straight Waveguide" sch_x=157 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16932 N$33863 N$33864 "Straight Waveguide" sch_x=157 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16933 N$33865 N$33866 "Straight Waveguide" sch_x=157 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16934 N$33867 N$33868 "Straight Waveguide" sch_x=157 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16935 N$33869 N$33870 "Straight Waveguide" sch_x=157 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16936 N$33871 N$33872 "Straight Waveguide" sch_x=157 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16937 N$33873 N$33874 "Straight Waveguide" sch_x=157 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16938 N$33875 N$33876 "Straight Waveguide" sch_x=157 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16939 N$33877 N$33878 "Straight Waveguide" sch_x=157 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16940 N$33879 N$33880 "Straight Waveguide" sch_x=157 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16941 N$33881 N$33882 "Straight Waveguide" sch_x=157 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16942 N$33883 N$33884 "Straight Waveguide" sch_x=157 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16943 N$33885 N$33886 "Straight Waveguide" sch_x=155 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16944 N$33887 N$33888 "Straight Waveguide" sch_x=155 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16945 N$33889 N$33890 "Straight Waveguide" sch_x=155 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16946 N$33891 N$33892 "Straight Waveguide" sch_x=155 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16947 N$33893 N$33894 "Straight Waveguide" sch_x=155 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16948 N$33895 N$33896 "Straight Waveguide" sch_x=155 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16949 N$33897 N$33898 "Straight Waveguide" sch_x=155 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16950 N$33899 N$33900 "Straight Waveguide" sch_x=155 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16951 N$33901 N$33902 "Straight Waveguide" sch_x=155 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16952 N$33903 N$33904 "Straight Waveguide" sch_x=155 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16953 N$33905 N$33906 "Straight Waveguide" sch_x=155 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16954 N$33907 N$33908 "Straight Waveguide" sch_x=155 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16955 N$33909 N$33910 "Straight Waveguide" sch_x=155 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16956 N$33911 N$33912 "Straight Waveguide" sch_x=155 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16957 N$33913 N$33914 "Straight Waveguide" sch_x=155 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16958 N$33915 N$33916 "Straight Waveguide" sch_x=155 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16959 N$33917 N$33918 "Straight Waveguide" sch_x=155 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16960 N$33919 N$33920 "Straight Waveguide" sch_x=155 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16961 N$33921 N$33922 "Straight Waveguide" sch_x=155 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16962 N$33923 N$33924 "Straight Waveguide" sch_x=155 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16963 N$33925 N$33926 "Straight Waveguide" sch_x=155 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16964 N$33927 N$33928 "Straight Waveguide" sch_x=155 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16965 N$33929 N$33930 "Straight Waveguide" sch_x=155 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16966 N$33931 N$33932 "Straight Waveguide" sch_x=155 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16967 N$33933 N$33934 "Straight Waveguide" sch_x=155 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16968 N$33935 N$33936 "Straight Waveguide" sch_x=155 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16969 N$33937 N$33938 "Straight Waveguide" sch_x=155 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16970 N$33939 N$33940 "Straight Waveguide" sch_x=155 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16971 N$33941 N$33942 "Straight Waveguide" sch_x=153 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16972 N$33943 N$33944 "Straight Waveguide" sch_x=153 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16973 N$33945 N$33946 "Straight Waveguide" sch_x=153 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16974 N$33947 N$33948 "Straight Waveguide" sch_x=153 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16975 N$33949 N$33950 "Straight Waveguide" sch_x=153 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16976 N$33951 N$33952 "Straight Waveguide" sch_x=153 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16977 N$33953 N$33954 "Straight Waveguide" sch_x=153 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16978 N$33955 N$33956 "Straight Waveguide" sch_x=153 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16979 N$33957 N$33958 "Straight Waveguide" sch_x=153 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16980 N$33959 N$33960 "Straight Waveguide" sch_x=153 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16981 N$33961 N$33962 "Straight Waveguide" sch_x=153 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16982 N$33963 N$33964 "Straight Waveguide" sch_x=153 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16983 N$33965 N$33966 "Straight Waveguide" sch_x=153 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16984 N$33967 N$33968 "Straight Waveguide" sch_x=153 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16985 N$33969 N$33970 "Straight Waveguide" sch_x=153 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16986 N$33971 N$33972 "Straight Waveguide" sch_x=153 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16987 N$33973 N$33974 "Straight Waveguide" sch_x=153 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16988 N$33975 N$33976 "Straight Waveguide" sch_x=153 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16989 N$33977 N$33978 "Straight Waveguide" sch_x=153 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16990 N$33979 N$33980 "Straight Waveguide" sch_x=153 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16991 N$33981 N$33982 "Straight Waveguide" sch_x=153 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16992 N$33983 N$33984 "Straight Waveguide" sch_x=153 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16993 N$33985 N$33986 "Straight Waveguide" sch_x=153 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16994 N$33987 N$33988 "Straight Waveguide" sch_x=153 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16995 N$33989 N$33990 "Straight Waveguide" sch_x=153 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16996 N$33991 N$33992 "Straight Waveguide" sch_x=153 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16997 N$33993 N$33994 "Straight Waveguide" sch_x=151 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16998 N$33995 N$33996 "Straight Waveguide" sch_x=151 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16999 N$33997 N$33998 "Straight Waveguide" sch_x=151 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17000 N$33999 N$34000 "Straight Waveguide" sch_x=151 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17001 N$34001 N$34002 "Straight Waveguide" sch_x=151 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17002 N$34003 N$34004 "Straight Waveguide" sch_x=151 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17003 N$34005 N$34006 "Straight Waveguide" sch_x=151 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17004 N$34007 N$34008 "Straight Waveguide" sch_x=151 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17005 N$34009 N$34010 "Straight Waveguide" sch_x=151 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17006 N$34011 N$34012 "Straight Waveguide" sch_x=151 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17007 N$34013 N$34014 "Straight Waveguide" sch_x=151 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17008 N$34015 N$34016 "Straight Waveguide" sch_x=151 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17009 N$34017 N$34018 "Straight Waveguide" sch_x=151 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17010 N$34019 N$34020 "Straight Waveguide" sch_x=151 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17011 N$34021 N$34022 "Straight Waveguide" sch_x=151 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17012 N$34023 N$34024 "Straight Waveguide" sch_x=151 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17013 N$34025 N$34026 "Straight Waveguide" sch_x=151 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17014 N$34027 N$34028 "Straight Waveguide" sch_x=151 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17015 N$34029 N$34030 "Straight Waveguide" sch_x=151 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17016 N$34031 N$34032 "Straight Waveguide" sch_x=151 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17017 N$34033 N$34034 "Straight Waveguide" sch_x=151 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17018 N$34035 N$34036 "Straight Waveguide" sch_x=151 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17019 N$34037 N$34038 "Straight Waveguide" sch_x=151 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17020 N$34039 N$34040 "Straight Waveguide" sch_x=151 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17021 N$34041 N$34042 "Straight Waveguide" sch_x=149 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17022 N$34043 N$34044 "Straight Waveguide" sch_x=149 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17023 N$34045 N$34046 "Straight Waveguide" sch_x=149 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17024 N$34047 N$34048 "Straight Waveguide" sch_x=149 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17025 N$34049 N$34050 "Straight Waveguide" sch_x=149 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17026 N$34051 N$34052 "Straight Waveguide" sch_x=149 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17027 N$34053 N$34054 "Straight Waveguide" sch_x=149 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17028 N$34055 N$34056 "Straight Waveguide" sch_x=149 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17029 N$34057 N$34058 "Straight Waveguide" sch_x=149 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17030 N$34059 N$34060 "Straight Waveguide" sch_x=149 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17031 N$34061 N$34062 "Straight Waveguide" sch_x=149 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17032 N$34063 N$34064 "Straight Waveguide" sch_x=149 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17033 N$34065 N$34066 "Straight Waveguide" sch_x=149 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17034 N$34067 N$34068 "Straight Waveguide" sch_x=149 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17035 N$34069 N$34070 "Straight Waveguide" sch_x=149 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17036 N$34071 N$34072 "Straight Waveguide" sch_x=149 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17037 N$34073 N$34074 "Straight Waveguide" sch_x=149 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17038 N$34075 N$34076 "Straight Waveguide" sch_x=149 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17039 N$34077 N$34078 "Straight Waveguide" sch_x=149 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17040 N$34079 N$34080 "Straight Waveguide" sch_x=149 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17041 N$34081 N$34082 "Straight Waveguide" sch_x=149 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17042 N$34083 N$34084 "Straight Waveguide" sch_x=149 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17043 N$34085 N$34086 "Straight Waveguide" sch_x=147 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17044 N$34087 N$34088 "Straight Waveguide" sch_x=147 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17045 N$34089 N$34090 "Straight Waveguide" sch_x=147 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17046 N$34091 N$34092 "Straight Waveguide" sch_x=147 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17047 N$34093 N$34094 "Straight Waveguide" sch_x=147 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17048 N$34095 N$34096 "Straight Waveguide" sch_x=147 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17049 N$34097 N$34098 "Straight Waveguide" sch_x=147 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17050 N$34099 N$34100 "Straight Waveguide" sch_x=147 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17051 N$34101 N$34102 "Straight Waveguide" sch_x=147 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17052 N$34103 N$34104 "Straight Waveguide" sch_x=147 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17053 N$34105 N$34106 "Straight Waveguide" sch_x=147 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17054 N$34107 N$34108 "Straight Waveguide" sch_x=147 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17055 N$34109 N$34110 "Straight Waveguide" sch_x=147 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17056 N$34111 N$34112 "Straight Waveguide" sch_x=147 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17057 N$34113 N$34114 "Straight Waveguide" sch_x=147 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17058 N$34115 N$34116 "Straight Waveguide" sch_x=147 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17059 N$34117 N$34118 "Straight Waveguide" sch_x=147 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17060 N$34119 N$34120 "Straight Waveguide" sch_x=147 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17061 N$34121 N$34122 "Straight Waveguide" sch_x=147 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17062 N$34123 N$34124 "Straight Waveguide" sch_x=147 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17063 N$34125 N$34126 "Straight Waveguide" sch_x=145 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17064 N$34127 N$34128 "Straight Waveguide" sch_x=145 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17065 N$34129 N$34130 "Straight Waveguide" sch_x=145 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17066 N$34131 N$34132 "Straight Waveguide" sch_x=145 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17067 N$34133 N$34134 "Straight Waveguide" sch_x=145 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17068 N$34135 N$34136 "Straight Waveguide" sch_x=145 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17069 N$34137 N$34138 "Straight Waveguide" sch_x=145 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17070 N$34139 N$34140 "Straight Waveguide" sch_x=145 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17071 N$34141 N$34142 "Straight Waveguide" sch_x=145 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17072 N$34143 N$34144 "Straight Waveguide" sch_x=145 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17073 N$34145 N$34146 "Straight Waveguide" sch_x=145 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17074 N$34147 N$34148 "Straight Waveguide" sch_x=145 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17075 N$34149 N$34150 "Straight Waveguide" sch_x=145 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17076 N$34151 N$34152 "Straight Waveguide" sch_x=145 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17077 N$34153 N$34154 "Straight Waveguide" sch_x=145 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17078 N$34155 N$34156 "Straight Waveguide" sch_x=145 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17079 N$34157 N$34158 "Straight Waveguide" sch_x=145 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17080 N$34159 N$34160 "Straight Waveguide" sch_x=145 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17081 N$34161 N$34162 "Straight Waveguide" sch_x=143 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17082 N$34163 N$34164 "Straight Waveguide" sch_x=143 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17083 N$34165 N$34166 "Straight Waveguide" sch_x=143 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17084 N$34167 N$34168 "Straight Waveguide" sch_x=143 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17085 N$34169 N$34170 "Straight Waveguide" sch_x=143 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17086 N$34171 N$34172 "Straight Waveguide" sch_x=143 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17087 N$34173 N$34174 "Straight Waveguide" sch_x=143 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17088 N$34175 N$34176 "Straight Waveguide" sch_x=143 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17089 N$34177 N$34178 "Straight Waveguide" sch_x=143 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17090 N$34179 N$34180 "Straight Waveguide" sch_x=143 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17091 N$34181 N$34182 "Straight Waveguide" sch_x=143 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17092 N$34183 N$34184 "Straight Waveguide" sch_x=143 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17093 N$34185 N$34186 "Straight Waveguide" sch_x=143 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17094 N$34187 N$34188 "Straight Waveguide" sch_x=143 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17095 N$34189 N$34190 "Straight Waveguide" sch_x=143 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17096 N$34191 N$34192 "Straight Waveguide" sch_x=143 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17097 N$34193 N$34194 "Straight Waveguide" sch_x=141 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17098 N$34195 N$34196 "Straight Waveguide" sch_x=141 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17099 N$34197 N$34198 "Straight Waveguide" sch_x=141 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17100 N$34199 N$34200 "Straight Waveguide" sch_x=141 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17101 N$34201 N$34202 "Straight Waveguide" sch_x=141 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17102 N$34203 N$34204 "Straight Waveguide" sch_x=141 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17103 N$34205 N$34206 "Straight Waveguide" sch_x=141 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17104 N$34207 N$34208 "Straight Waveguide" sch_x=141 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17105 N$34209 N$34210 "Straight Waveguide" sch_x=141 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17106 N$34211 N$34212 "Straight Waveguide" sch_x=141 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17107 N$34213 N$34214 "Straight Waveguide" sch_x=141 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17108 N$34215 N$34216 "Straight Waveguide" sch_x=141 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17109 N$34217 N$34218 "Straight Waveguide" sch_x=141 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17110 N$34219 N$34220 "Straight Waveguide" sch_x=141 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17111 N$34221 N$34222 "Straight Waveguide" sch_x=139 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17112 N$34223 N$34224 "Straight Waveguide" sch_x=139 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17113 N$34225 N$34226 "Straight Waveguide" sch_x=139 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17114 N$34227 N$34228 "Straight Waveguide" sch_x=139 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17115 N$34229 N$34230 "Straight Waveguide" sch_x=139 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17116 N$34231 N$34232 "Straight Waveguide" sch_x=139 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17117 N$34233 N$34234 "Straight Waveguide" sch_x=139 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17118 N$34235 N$34236 "Straight Waveguide" sch_x=139 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17119 N$34237 N$34238 "Straight Waveguide" sch_x=139 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17120 N$34239 N$34240 "Straight Waveguide" sch_x=139 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17121 N$34241 N$34242 "Straight Waveguide" sch_x=139 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17122 N$34243 N$34244 "Straight Waveguide" sch_x=139 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17123 N$34245 N$34246 "Straight Waveguide" sch_x=137 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17124 N$34247 N$34248 "Straight Waveguide" sch_x=137 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17125 N$34249 N$34250 "Straight Waveguide" sch_x=137 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17126 N$34251 N$34252 "Straight Waveguide" sch_x=137 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17127 N$34253 N$34254 "Straight Waveguide" sch_x=137 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17128 N$34255 N$34256 "Straight Waveguide" sch_x=137 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17129 N$34257 N$34258 "Straight Waveguide" sch_x=137 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17130 N$34259 N$34260 "Straight Waveguide" sch_x=137 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17131 N$34261 N$34262 "Straight Waveguide" sch_x=137 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17132 N$34263 N$34264 "Straight Waveguide" sch_x=137 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17133 N$34265 N$34266 "Straight Waveguide" sch_x=135 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17134 N$34267 N$34268 "Straight Waveguide" sch_x=135 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17135 N$34269 N$34270 "Straight Waveguide" sch_x=135 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17136 N$34271 N$34272 "Straight Waveguide" sch_x=135 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17137 N$34273 N$34274 "Straight Waveguide" sch_x=135 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17138 N$34275 N$34276 "Straight Waveguide" sch_x=135 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17139 N$34277 N$34278 "Straight Waveguide" sch_x=135 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17140 N$34279 N$34280 "Straight Waveguide" sch_x=135 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17141 N$34281 N$34282 "Straight Waveguide" sch_x=133 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17142 N$34283 N$34284 "Straight Waveguide" sch_x=133 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17143 N$34285 N$34286 "Straight Waveguide" sch_x=133 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17144 N$34287 N$34288 "Straight Waveguide" sch_x=133 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17145 N$34289 N$34290 "Straight Waveguide" sch_x=133 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17146 N$34291 N$34292 "Straight Waveguide" sch_x=133 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17147 N$34293 N$34294 "Straight Waveguide" sch_x=131 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17148 N$34295 N$34296 "Straight Waveguide" sch_x=131 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17149 N$34297 N$34298 "Straight Waveguide" sch_x=131 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17150 N$34299 N$34300 "Straight Waveguide" sch_x=131 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17151 N$34301 N$34302 "Straight Waveguide" sch_x=129 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17152 N$34303 N$34304 "Straight Waveguide" sch_x=129 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17153 N$34306 N$34305 "Straight Waveguide" sch_x=189 sch_y=62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17154 N$34308 N$34307 "Straight Waveguide" sch_x=188 sch_y=61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17155 N$34310 N$34309 "Straight Waveguide" sch_x=187 sch_y=60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17156 N$34312 N$34311 "Straight Waveguide" sch_x=186 sch_y=59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17157 N$34314 N$34313 "Straight Waveguide" sch_x=185 sch_y=58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17158 N$34316 N$34315 "Straight Waveguide" sch_x=184 sch_y=57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17159 N$34318 N$34317 "Straight Waveguide" sch_x=183 sch_y=56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17160 N$34320 N$34319 "Straight Waveguide" sch_x=182 sch_y=55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17161 N$34322 N$34321 "Straight Waveguide" sch_x=181 sch_y=54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17162 N$34324 N$34323 "Straight Waveguide" sch_x=180 sch_y=53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17163 N$34326 N$34325 "Straight Waveguide" sch_x=179 sch_y=52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17164 N$34328 N$34327 "Straight Waveguide" sch_x=178 sch_y=51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17165 N$34330 N$34329 "Straight Waveguide" sch_x=177 sch_y=50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17166 N$34332 N$34331 "Straight Waveguide" sch_x=176 sch_y=49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17167 N$34334 N$34333 "Straight Waveguide" sch_x=175 sch_y=48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17168 N$34336 N$34335 "Straight Waveguide" sch_x=174 sch_y=47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17169 N$34338 N$34337 "Straight Waveguide" sch_x=173 sch_y=46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17170 N$34340 N$34339 "Straight Waveguide" sch_x=172 sch_y=45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17171 N$34342 N$34341 "Straight Waveguide" sch_x=171 sch_y=44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17172 N$34344 N$34343 "Straight Waveguide" sch_x=170 sch_y=43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17173 N$34346 N$34345 "Straight Waveguide" sch_x=169 sch_y=42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17174 N$34348 N$34347 "Straight Waveguide" sch_x=168 sch_y=41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17175 N$34350 N$34349 "Straight Waveguide" sch_x=167 sch_y=40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17176 N$34352 N$34351 "Straight Waveguide" sch_x=166 sch_y=39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17177 N$34354 N$34353 "Straight Waveguide" sch_x=165 sch_y=38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17178 N$34356 N$34355 "Straight Waveguide" sch_x=164 sch_y=37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17179 N$34358 N$34357 "Straight Waveguide" sch_x=163 sch_y=36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17180 N$34360 N$34359 "Straight Waveguide" sch_x=162 sch_y=35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17181 N$34362 N$34361 "Straight Waveguide" sch_x=161 sch_y=34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17182 N$34364 N$34363 "Straight Waveguide" sch_x=160 sch_y=33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17183 N$34366 N$34365 "Straight Waveguide" sch_x=159 sch_y=32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17184 N$34368 N$34367 "Straight Waveguide" sch_x=158 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17185 N$34370 N$34369 "Straight Waveguide" sch_x=157 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17186 N$34372 N$34371 "Straight Waveguide" sch_x=156 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17187 N$34374 N$34373 "Straight Waveguide" sch_x=155 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17188 N$34376 N$34375 "Straight Waveguide" sch_x=154 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17189 N$34378 N$34377 "Straight Waveguide" sch_x=153 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17190 N$34380 N$34379 "Straight Waveguide" sch_x=152 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17191 N$34382 N$34381 "Straight Waveguide" sch_x=151 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17192 N$34384 N$34383 "Straight Waveguide" sch_x=150 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17193 N$34386 N$34385 "Straight Waveguide" sch_x=149 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17194 N$34388 N$34387 "Straight Waveguide" sch_x=148 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17195 N$34390 N$34389 "Straight Waveguide" sch_x=147 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17196 N$34392 N$34391 "Straight Waveguide" sch_x=146 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17197 N$34394 N$34393 "Straight Waveguide" sch_x=145 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17198 N$34396 N$34395 "Straight Waveguide" sch_x=144 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17199 N$34398 N$34397 "Straight Waveguide" sch_x=143 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17200 N$34400 N$34399 "Straight Waveguide" sch_x=142 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17201 N$34402 N$34401 "Straight Waveguide" sch_x=141 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17202 N$34404 N$34403 "Straight Waveguide" sch_x=140 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17203 N$34406 N$34405 "Straight Waveguide" sch_x=139 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17204 N$34408 N$34407 "Straight Waveguide" sch_x=138 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17205 N$34410 N$34409 "Straight Waveguide" sch_x=137 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17206 N$34412 N$34411 "Straight Waveguide" sch_x=136 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17207 N$34414 N$34413 "Straight Waveguide" sch_x=135 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17208 N$34416 N$34415 "Straight Waveguide" sch_x=134 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17209 N$34418 N$34417 "Straight Waveguide" sch_x=133 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17210 N$34420 N$34419 "Straight Waveguide" sch_x=132 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17211 N$34422 N$34421 "Straight Waveguide" sch_x=131 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17212 N$34424 N$34423 "Straight Waveguide" sch_x=130 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17213 N$34426 N$34425 "Straight Waveguide" sch_x=129 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17214 N$34428 N$34427 "Straight Waveguide" sch_x=128 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17215 N$34430 N$34429 "Straight Waveguide" sch_x=127 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17216 N$34432 N$34431 "Straight Waveguide" sch_x=127 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17217 N$34434 N$34433 "Straight Waveguide" sch_x=128 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17218 N$34436 N$34435 "Straight Waveguide" sch_x=129 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17219 N$34438 N$34437 "Straight Waveguide" sch_x=130 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17220 N$34440 N$34439 "Straight Waveguide" sch_x=131 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17221 N$34442 N$34441 "Straight Waveguide" sch_x=132 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17222 N$34444 N$34443 "Straight Waveguide" sch_x=133 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17223 N$34446 N$34445 "Straight Waveguide" sch_x=134 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17224 N$34448 N$34447 "Straight Waveguide" sch_x=135 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17225 N$34450 N$34449 "Straight Waveguide" sch_x=136 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17226 N$34452 N$34451 "Straight Waveguide" sch_x=137 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17227 N$34454 N$34453 "Straight Waveguide" sch_x=138 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17228 N$34456 N$34455 "Straight Waveguide" sch_x=139 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17229 N$34458 N$34457 "Straight Waveguide" sch_x=140 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17230 N$34460 N$34459 "Straight Waveguide" sch_x=141 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17231 N$34462 N$34461 "Straight Waveguide" sch_x=142 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17232 N$34464 N$34463 "Straight Waveguide" sch_x=143 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17233 N$34466 N$34465 "Straight Waveguide" sch_x=144 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17234 N$34468 N$34467 "Straight Waveguide" sch_x=145 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17235 N$34470 N$34469 "Straight Waveguide" sch_x=146 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17236 N$34472 N$34471 "Straight Waveguide" sch_x=147 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17237 N$34474 N$34473 "Straight Waveguide" sch_x=148 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17238 N$34476 N$34475 "Straight Waveguide" sch_x=149 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17239 N$34478 N$34477 "Straight Waveguide" sch_x=150 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17240 N$34480 N$34479 "Straight Waveguide" sch_x=151 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17241 N$34482 N$34481 "Straight Waveguide" sch_x=152 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17242 N$34484 N$34483 "Straight Waveguide" sch_x=153 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17243 N$34486 N$34485 "Straight Waveguide" sch_x=154 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17244 N$34488 N$34487 "Straight Waveguide" sch_x=155 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17245 N$34490 N$34489 "Straight Waveguide" sch_x=156 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17246 N$34492 N$34491 "Straight Waveguide" sch_x=157 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17247 N$34494 N$34493 "Straight Waveguide" sch_x=158 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17248 N$34496 N$34495 "Straight Waveguide" sch_x=159 sch_y=-32.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17249 N$34498 N$34497 "Straight Waveguide" sch_x=160 sch_y=-33 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17250 N$34500 N$34499 "Straight Waveguide" sch_x=161 sch_y=-34.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17251 N$34502 N$34501 "Straight Waveguide" sch_x=162 sch_y=-35 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17252 N$34504 N$34503 "Straight Waveguide" sch_x=163 sch_y=-36.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17253 N$34506 N$34505 "Straight Waveguide" sch_x=164 sch_y=-37 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17254 N$34508 N$34507 "Straight Waveguide" sch_x=165 sch_y=-38.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17255 N$34510 N$34509 "Straight Waveguide" sch_x=166 sch_y=-39 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17256 N$34512 N$34511 "Straight Waveguide" sch_x=167 sch_y=-40.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17257 N$34514 N$34513 "Straight Waveguide" sch_x=168 sch_y=-41 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17258 N$34516 N$34515 "Straight Waveguide" sch_x=169 sch_y=-42.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17259 N$34518 N$34517 "Straight Waveguide" sch_x=170 sch_y=-43 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17260 N$34520 N$34519 "Straight Waveguide" sch_x=171 sch_y=-44.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17261 N$34522 N$34521 "Straight Waveguide" sch_x=172 sch_y=-45 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17262 N$34524 N$34523 "Straight Waveguide" sch_x=173 sch_y=-46.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17263 N$34526 N$34525 "Straight Waveguide" sch_x=174 sch_y=-47 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17264 N$34528 N$34527 "Straight Waveguide" sch_x=175 sch_y=-48.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17265 N$34530 N$34529 "Straight Waveguide" sch_x=176 sch_y=-49 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17266 N$34532 N$34531 "Straight Waveguide" sch_x=177 sch_y=-50.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17267 N$34534 N$34533 "Straight Waveguide" sch_x=178 sch_y=-51 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17268 N$34536 N$34535 "Straight Waveguide" sch_x=179 sch_y=-52.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17269 N$34538 N$34537 "Straight Waveguide" sch_x=180 sch_y=-53 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17270 N$34540 N$34539 "Straight Waveguide" sch_x=181 sch_y=-54.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17271 N$34542 N$34541 "Straight Waveguide" sch_x=182 sch_y=-55 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17272 N$34544 N$34543 "Straight Waveguide" sch_x=183 sch_y=-56.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17273 N$34546 N$34545 "Straight Waveguide" sch_x=184 sch_y=-57 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17274 N$34548 N$34547 "Straight Waveguide" sch_x=185 sch_y=-58.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17275 N$34550 N$34549 "Straight Waveguide" sch_x=186 sch_y=-59 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17276 N$34552 N$34551 "Straight Waveguide" sch_x=187 sch_y=-60.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17277 N$34554 N$34553 "Straight Waveguide" sch_x=188 sch_y=-61 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17278 N$34556 N$34555 "Straight Waveguide" sch_x=189 sch_y=-62.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17279 N$34558 N$34557 "Straight Waveguide" sch_x=190 sch_y=63 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17280 N$34560 N$34559 "Straight Waveguide" sch_x=190 sch_y=-63 sch_r=0 sch_f=false lay_x=0 lay_y=0
.ends HDBE
* - ONA
.ona input_unit=wavelength input_parameter=center_and_range center=1550e-9
  + range=100e-9 number_of_points=100 
  + minimum_loss=200
  + sensitivity=-200 
  + analysis_type=scattering_data
  + multithreading=user_defined number_of_threads=1 
 + input(1)=HDBE,N$34945
+ input(2)=HDBE,N$34947
+ input(3)=HDBE,N$34949
+ input(4)=HDBE,N$34951
+ input(5)=HDBE,N$34953
+ input(6)=HDBE,N$34955
+ input(7)=HDBE,N$34957
+ input(8)=HDBE,N$34959
+ input(9)=HDBE,N$34961
+ input(10)=HDBE,N$34963
+ input(11)=HDBE,N$34965
+ input(12)=HDBE,N$34967
+ input(13)=HDBE,N$34969
+ input(14)=HDBE,N$34971
+ input(15)=HDBE,N$34973
+ input(16)=HDBE,N$34975
+ input(17)=HDBE,N$34977
+ input(18)=HDBE,N$34979
+ input(19)=HDBE,N$34981
+ input(20)=HDBE,N$34983
+ input(21)=HDBE,N$34985
+ input(22)=HDBE,N$34987
+ input(23)=HDBE,N$34989
+ input(24)=HDBE,N$34991
+ input(25)=HDBE,N$34993
+ input(26)=HDBE,N$34995
+ input(27)=HDBE,N$34997
+ input(28)=HDBE,N$34999
+ input(29)=HDBE,N$35001
+ input(30)=HDBE,N$35003
+ input(31)=HDBE,N$35005
+ input(32)=HDBE,N$35007
+ input(33)=HDBE,N$35009
+ input(34)=HDBE,N$35011
+ input(35)=HDBE,N$35013
+ input(36)=HDBE,N$35015
+ input(37)=HDBE,N$35017
+ input(38)=HDBE,N$35019
+ input(39)=HDBE,N$35021
+ input(40)=HDBE,N$35023
+ input(41)=HDBE,N$35025
+ input(42)=HDBE,N$35027
+ input(43)=HDBE,N$35029
+ input(44)=HDBE,N$35031
+ input(45)=HDBE,N$35033
+ input(46)=HDBE,N$35035
+ input(47)=HDBE,N$35037
+ input(48)=HDBE,N$35039
+ input(49)=HDBE,N$35041
+ input(50)=HDBE,N$35043
+ input(51)=HDBE,N$35045
+ input(52)=HDBE,N$35047
+ input(53)=HDBE,N$35049
+ input(54)=HDBE,N$35051
+ input(55)=HDBE,N$35053
+ input(56)=HDBE,N$35055
+ input(57)=HDBE,N$35057
+ input(58)=HDBE,N$35059
+ input(59)=HDBE,N$35061
+ input(60)=HDBE,N$35063
+ input(61)=HDBE,N$35065
+ input(62)=HDBE,N$35067
+ input(63)=HDBE,N$35069
+ input(64)=HDBE,N$35071
  + output=HDBE,N$34561

HDBE  N$34561 N$34563 N$34565 N$34567 N$34569 N$34571 N$34573 N$34575 N$34577 N$34579 N$34581 N$34583 N$34585 N$34587 N$34589 N$34591 N$34593 N$34595 N$34597 N$34599 N$34601 N$34603 N$34605 N$34607 N$34609 N$34611 N$34613 N$34615 N$34617 N$34619 N$34621 N$34623 N$34625 N$34627 N$34629 N$34631 N$34633 N$34635 N$34637 N$34639 N$34641 N$34643 N$34645 N$34647 N$34649 N$34651 N$34653 N$34655 N$34657 N$34659 N$34661 N$34663 N$34665 N$34667 N$34669 N$34671 N$34673 N$34675 N$34677 N$34679 N$34681 N$34683 N$34685 N$34687 N$34945 N$34947 N$34949 N$34951 N$34953 N$34955 N$34957 N$34959 N$34961 N$34963 N$34965 N$34967 N$34969 N$34971 N$34973 N$34975 N$34977 N$34979 N$34981 N$34983 N$34985 N$34987 N$34989 N$34991 N$34993 N$34995 N$34997 N$34999 N$35001 N$35003 N$35005 N$35007 N$35009 N$35011 N$35013 N$35015 N$35017 N$35019 N$35021 N$35023 N$35025 N$35027 N$35029 N$35031 N$35033 N$35035 N$35037 N$35039 N$35041 N$35043 N$35045 N$35047 N$35049 N$35051 N$35053 N$35055 N$35057 N$35059 N$35061 N$35063 N$35065 N$35067 N$35069 N$35071 HDBE sch_x=0 sch_y=0
*
.end