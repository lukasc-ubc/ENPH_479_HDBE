*
* MAIN CELL: Component pathname : root_element
*
   .MODEL BDC_switch_ideal "label 1"="TE" "control"=1
   .MODEL "Waveguide Crossing" "label 1"="TE" "transmission 1"=0.9954054174 "cross talk 1"=0.0001
   + "transmission 2"=1 "cross talk 2"=0 "reflection 1"=0.001
   + "reflection 2"=0 "label 2"="TM" "orthogonal identifier 1"=1
   + "orthogonal identifier 2"=2
   .MODEL "Straight Waveguide" "excess loss temperature sensitivity 2"=0 "label 1"="TE" "orthogonal identifier 1"=1 
   + "loss 1"=0 "number of taps"=64 "dispersion 1"=0 
   + "effective index temperature sensitivity 2"=0 "effective index 2"=1 length=10u 
   + "group index 2"=1 "orthogonal identifier 2"=2 "nominal temperature"=300 
   + "loss 2"=0 "dispersion 2"=0 frequency=193.1T 
   + "digital filter"=0 "run diagnostic"=0 "window function"="rectangular" 
   + "thermal fill factor"=1 "excess loss temperature sensitivity 1"=0 "label 2"="TM" 
   + "thermal effects"=0 "effective index temperature sensitivity 1"=0 "effective index 1"=1 

.subckt HDBE  N$2369 N$2371 N$2373 N$2375 N$2377 N$2379 N$2381 N$2383 N$2385 N$2387 N$2389 N$2391 N$2393 N$2395 N$2397 N$2399 N$2465 N$2467 N$2469 N$2471 N$2473 N$2475 N$2477 N$2479 N$2481 N$2483 N$2485 N$2487 N$2489 N$2491 N$2493 N$2495
   S353 N$2369 N$2370 N$1821 N$1282 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S354 N$2371 N$2372 N$1284 N$1286 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S355 N$2373 N$2374 N$1288 N$1290 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S356 N$2375 N$2376 N$1292 N$1294 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S357 N$2377 N$2378 N$1296 N$1298 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S358 N$2379 N$2380 N$1300 N$1302 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S359 N$2381 N$2382 N$1304 N$1306 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S360 N$2383 N$2384 N$1308 N$1310 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S361 N$2385 N$2386 N$1312 N$1314 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S362 N$2387 N$2388 N$1316 N$1318 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S363 N$2389 N$2390 N$1320 N$1322 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S364 N$2391 N$2392 N$1324 N$1326 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S365 N$2393 N$2394 N$1328 N$1330 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S366 N$2395 N$2396 N$1332 N$1334 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S367 N$2397 N$2398 N$1336 N$1338 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S368 N$2399 N$2400 N$1340 N$1823 BDC_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C369 N$1281 N$1283 N$1761 N$1342 "Waveguide Crossing" sch_x=-60 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C370 N$1285 N$1287 N$1344 N$1346 "Waveguide Crossing" sch_x=-60 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C371 N$1289 N$1291 N$1348 N$1350 "Waveguide Crossing" sch_x=-60 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C372 N$1293 N$1295 N$1352 N$1354 "Waveguide Crossing" sch_x=-60 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C373 N$1297 N$1299 N$1356 N$1358 "Waveguide Crossing" sch_x=-60 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C374 N$1301 N$1303 N$1360 N$1362 "Waveguide Crossing" sch_x=-60 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C375 N$1305 N$1307 N$1364 N$1366 "Waveguide Crossing" sch_x=-60 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C376 N$1309 N$1311 N$1368 N$1370 "Waveguide Crossing" sch_x=-60 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C377 N$1313 N$1315 N$1372 N$1374 "Waveguide Crossing" sch_x=-60 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C378 N$1317 N$1319 N$1376 N$1378 "Waveguide Crossing" sch_x=-60 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C379 N$1321 N$1323 N$1380 N$1382 "Waveguide Crossing" sch_x=-60 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C380 N$1325 N$1327 N$1384 N$1386 "Waveguide Crossing" sch_x=-60 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C381 N$1329 N$1331 N$1388 N$1390 "Waveguide Crossing" sch_x=-60 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C382 N$1333 N$1335 N$1392 N$1394 "Waveguide Crossing" sch_x=-60 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C383 N$1337 N$1339 N$1396 N$1819 "Waveguide Crossing" sch_x=-60 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C384 N$1341 N$1343 N$1763 N$1398 "Waveguide Crossing" sch_x=-58 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C385 N$1345 N$1347 N$1400 N$1402 "Waveguide Crossing" sch_x=-58 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C386 N$1349 N$1351 N$1404 N$1406 "Waveguide Crossing" sch_x=-58 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C387 N$1353 N$1355 N$1408 N$1410 "Waveguide Crossing" sch_x=-58 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C388 N$1357 N$1359 N$1412 N$1414 "Waveguide Crossing" sch_x=-58 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C389 N$1361 N$1363 N$1416 N$1418 "Waveguide Crossing" sch_x=-58 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C390 N$1365 N$1367 N$1420 N$1422 "Waveguide Crossing" sch_x=-58 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C391 N$1369 N$1371 N$1424 N$1426 "Waveguide Crossing" sch_x=-58 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C392 N$1373 N$1375 N$1428 N$1430 "Waveguide Crossing" sch_x=-58 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C393 N$1377 N$1379 N$1432 N$1434 "Waveguide Crossing" sch_x=-58 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C394 N$1381 N$1383 N$1436 N$1438 "Waveguide Crossing" sch_x=-58 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C395 N$1385 N$1387 N$1440 N$1442 "Waveguide Crossing" sch_x=-58 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C396 N$1389 N$1391 N$1444 N$1446 "Waveguide Crossing" sch_x=-58 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C397 N$1393 N$1395 N$1448 N$1817 "Waveguide Crossing" sch_x=-58 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C398 N$1397 N$1399 N$1765 N$1450 "Waveguide Crossing" sch_x=-56 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C399 N$1401 N$1403 N$1452 N$1454 "Waveguide Crossing" sch_x=-56 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C400 N$1405 N$1407 N$1456 N$1458 "Waveguide Crossing" sch_x=-56 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C401 N$1409 N$1411 N$1460 N$1462 "Waveguide Crossing" sch_x=-56 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C402 N$1413 N$1415 N$1464 N$1466 "Waveguide Crossing" sch_x=-56 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C403 N$1417 N$1419 N$1468 N$1470 "Waveguide Crossing" sch_x=-56 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C404 N$1421 N$1423 N$1472 N$1474 "Waveguide Crossing" sch_x=-56 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C405 N$1425 N$1427 N$1476 N$1478 "Waveguide Crossing" sch_x=-56 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C406 N$1429 N$1431 N$1480 N$1482 "Waveguide Crossing" sch_x=-56 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C407 N$1433 N$1435 N$1484 N$1486 "Waveguide Crossing" sch_x=-56 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C408 N$1437 N$1439 N$1488 N$1490 "Waveguide Crossing" sch_x=-56 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C409 N$1441 N$1443 N$1492 N$1494 "Waveguide Crossing" sch_x=-56 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C410 N$1445 N$1447 N$1496 N$1815 "Waveguide Crossing" sch_x=-56 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C411 N$1449 N$1451 N$1767 N$1498 "Waveguide Crossing" sch_x=-54 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C412 N$1453 N$1455 N$1500 N$1502 "Waveguide Crossing" sch_x=-54 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C413 N$1457 N$1459 N$1504 N$1506 "Waveguide Crossing" sch_x=-54 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C414 N$1461 N$1463 N$1508 N$1510 "Waveguide Crossing" sch_x=-54 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C415 N$1465 N$1467 N$1512 N$1514 "Waveguide Crossing" sch_x=-54 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C416 N$1469 N$1471 N$1516 N$1518 "Waveguide Crossing" sch_x=-54 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C417 N$1473 N$1475 N$1520 N$1522 "Waveguide Crossing" sch_x=-54 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C418 N$1477 N$1479 N$1524 N$1526 "Waveguide Crossing" sch_x=-54 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C419 N$1481 N$1483 N$1528 N$1530 "Waveguide Crossing" sch_x=-54 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C420 N$1485 N$1487 N$1532 N$1534 "Waveguide Crossing" sch_x=-54 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C421 N$1489 N$1491 N$1536 N$1538 "Waveguide Crossing" sch_x=-54 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C422 N$1493 N$1495 N$1540 N$1813 "Waveguide Crossing" sch_x=-54 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C423 N$1497 N$1499 N$1769 N$1542 "Waveguide Crossing" sch_x=-52 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C424 N$1501 N$1503 N$1544 N$1546 "Waveguide Crossing" sch_x=-52 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C425 N$1505 N$1507 N$1548 N$1550 "Waveguide Crossing" sch_x=-52 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C426 N$1509 N$1511 N$1552 N$1554 "Waveguide Crossing" sch_x=-52 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C427 N$1513 N$1515 N$1556 N$1558 "Waveguide Crossing" sch_x=-52 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C428 N$1517 N$1519 N$1560 N$1562 "Waveguide Crossing" sch_x=-52 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C429 N$1521 N$1523 N$1564 N$1566 "Waveguide Crossing" sch_x=-52 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C430 N$1525 N$1527 N$1568 N$1570 "Waveguide Crossing" sch_x=-52 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C431 N$1529 N$1531 N$1572 N$1574 "Waveguide Crossing" sch_x=-52 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C432 N$1533 N$1535 N$1576 N$1578 "Waveguide Crossing" sch_x=-52 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C433 N$1537 N$1539 N$1580 N$1811 "Waveguide Crossing" sch_x=-52 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C434 N$1541 N$1543 N$1771 N$1582 "Waveguide Crossing" sch_x=-50 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C435 N$1545 N$1547 N$1584 N$1586 "Waveguide Crossing" sch_x=-50 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C436 N$1549 N$1551 N$1588 N$1590 "Waveguide Crossing" sch_x=-50 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C437 N$1553 N$1555 N$1592 N$1594 "Waveguide Crossing" sch_x=-50 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C438 N$1557 N$1559 N$1596 N$1598 "Waveguide Crossing" sch_x=-50 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C439 N$1561 N$1563 N$1600 N$1602 "Waveguide Crossing" sch_x=-50 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C440 N$1565 N$1567 N$1604 N$1606 "Waveguide Crossing" sch_x=-50 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C441 N$1569 N$1571 N$1608 N$1610 "Waveguide Crossing" sch_x=-50 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C442 N$1573 N$1575 N$1612 N$1614 "Waveguide Crossing" sch_x=-50 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C443 N$1577 N$1579 N$1616 N$1809 "Waveguide Crossing" sch_x=-50 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C444 N$1581 N$1583 N$1773 N$1618 "Waveguide Crossing" sch_x=-48 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C445 N$1585 N$1587 N$1620 N$1622 "Waveguide Crossing" sch_x=-48 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C446 N$1589 N$1591 N$1624 N$1626 "Waveguide Crossing" sch_x=-48 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C447 N$1593 N$1595 N$1628 N$1630 "Waveguide Crossing" sch_x=-48 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C448 N$1597 N$1599 N$1632 N$1634 "Waveguide Crossing" sch_x=-48 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C449 N$1601 N$1603 N$1636 N$1638 "Waveguide Crossing" sch_x=-48 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C450 N$1605 N$1607 N$1640 N$1642 "Waveguide Crossing" sch_x=-48 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C451 N$1609 N$1611 N$1644 N$1646 "Waveguide Crossing" sch_x=-48 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C452 N$1613 N$1615 N$1648 N$1807 "Waveguide Crossing" sch_x=-48 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C453 N$1617 N$1619 N$1775 N$1650 "Waveguide Crossing" sch_x=-46 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C454 N$1621 N$1623 N$1652 N$1654 "Waveguide Crossing" sch_x=-46 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C455 N$1625 N$1627 N$1656 N$1658 "Waveguide Crossing" sch_x=-46 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C456 N$1629 N$1631 N$1660 N$1662 "Waveguide Crossing" sch_x=-46 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C457 N$1633 N$1635 N$1664 N$1666 "Waveguide Crossing" sch_x=-46 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C458 N$1637 N$1639 N$1668 N$1670 "Waveguide Crossing" sch_x=-46 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C459 N$1641 N$1643 N$1672 N$1674 "Waveguide Crossing" sch_x=-46 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C460 N$1645 N$1647 N$1676 N$1805 "Waveguide Crossing" sch_x=-46 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C461 N$1649 N$1651 N$1777 N$1678 "Waveguide Crossing" sch_x=-44 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C462 N$1653 N$1655 N$1680 N$1682 "Waveguide Crossing" sch_x=-44 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C463 N$1657 N$1659 N$1684 N$1686 "Waveguide Crossing" sch_x=-44 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C464 N$1661 N$1663 N$1688 N$1690 "Waveguide Crossing" sch_x=-44 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C465 N$1665 N$1667 N$1692 N$1694 "Waveguide Crossing" sch_x=-44 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C466 N$1669 N$1671 N$1696 N$1698 "Waveguide Crossing" sch_x=-44 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C467 N$1673 N$1675 N$1700 N$1803 "Waveguide Crossing" sch_x=-44 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C468 N$1677 N$1679 N$1779 N$1702 "Waveguide Crossing" sch_x=-42 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C469 N$1681 N$1683 N$1704 N$1706 "Waveguide Crossing" sch_x=-42 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C470 N$1685 N$1687 N$1708 N$1710 "Waveguide Crossing" sch_x=-42 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C471 N$1689 N$1691 N$1712 N$1714 "Waveguide Crossing" sch_x=-42 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C472 N$1693 N$1695 N$1716 N$1718 "Waveguide Crossing" sch_x=-42 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C473 N$1697 N$1699 N$1720 N$1801 "Waveguide Crossing" sch_x=-42 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C474 N$1701 N$1703 N$1781 N$1722 "Waveguide Crossing" sch_x=-40 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C475 N$1705 N$1707 N$1724 N$1726 "Waveguide Crossing" sch_x=-40 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C476 N$1709 N$1711 N$1728 N$1730 "Waveguide Crossing" sch_x=-40 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C477 N$1713 N$1715 N$1732 N$1734 "Waveguide Crossing" sch_x=-40 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C478 N$1717 N$1719 N$1736 N$1799 "Waveguide Crossing" sch_x=-40 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C479 N$1721 N$1723 N$1783 N$1738 "Waveguide Crossing" sch_x=-38 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C480 N$1725 N$1727 N$1740 N$1742 "Waveguide Crossing" sch_x=-38 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C481 N$1729 N$1731 N$1744 N$1746 "Waveguide Crossing" sch_x=-38 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C482 N$1733 N$1735 N$1748 N$1797 "Waveguide Crossing" sch_x=-38 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C483 N$1737 N$1739 N$1785 N$1750 "Waveguide Crossing" sch_x=-36 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C484 N$1741 N$1743 N$1752 N$1754 "Waveguide Crossing" sch_x=-36 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C485 N$1745 N$1747 N$1756 N$1795 "Waveguide Crossing" sch_x=-36 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C486 N$1749 N$1751 N$1787 N$1758 "Waveguide Crossing" sch_x=-34 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C487 N$1753 N$1755 N$1760 N$1793 "Waveguide Crossing" sch_x=-34 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C488 N$1757 N$1759 N$1789 N$1791 "Waveguide Crossing" sch_x=-32 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S281 N$1792 N$1794 N$1133 N$994 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S282 N$1796 N$1798 N$996 N$998 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S283 N$1800 N$1802 N$1000 N$1002 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S284 N$1804 N$1806 N$1004 N$1006 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S285 N$1808 N$1810 N$1008 N$1010 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S286 N$1812 N$1814 N$1012 N$1014 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S287 N$1816 N$1818 N$1016 N$1018 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S288 N$1820 N$1824 N$1020 N$1135 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C289 N$993 N$995 N$1105 N$1022 "Waveguide Crossing" sch_x=-28 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C290 N$997 N$999 N$1024 N$1026 "Waveguide Crossing" sch_x=-28 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C291 N$1001 N$1003 N$1028 N$1030 "Waveguide Crossing" sch_x=-28 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C292 N$1005 N$1007 N$1032 N$1034 "Waveguide Crossing" sch_x=-28 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C293 N$1009 N$1011 N$1036 N$1038 "Waveguide Crossing" sch_x=-28 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C294 N$1013 N$1015 N$1040 N$1042 "Waveguide Crossing" sch_x=-28 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C295 N$1017 N$1019 N$1044 N$1131 "Waveguide Crossing" sch_x=-28 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C296 N$1021 N$1023 N$1107 N$1046 "Waveguide Crossing" sch_x=-26 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C297 N$1025 N$1027 N$1048 N$1050 "Waveguide Crossing" sch_x=-26 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C298 N$1029 N$1031 N$1052 N$1054 "Waveguide Crossing" sch_x=-26 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C299 N$1033 N$1035 N$1056 N$1058 "Waveguide Crossing" sch_x=-26 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C300 N$1037 N$1039 N$1060 N$1062 "Waveguide Crossing" sch_x=-26 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C301 N$1041 N$1043 N$1064 N$1129 "Waveguide Crossing" sch_x=-26 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C302 N$1045 N$1047 N$1109 N$1066 "Waveguide Crossing" sch_x=-24 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C303 N$1049 N$1051 N$1068 N$1070 "Waveguide Crossing" sch_x=-24 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C304 N$1053 N$1055 N$1072 N$1074 "Waveguide Crossing" sch_x=-24 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C305 N$1057 N$1059 N$1076 N$1078 "Waveguide Crossing" sch_x=-24 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C306 N$1061 N$1063 N$1080 N$1127 "Waveguide Crossing" sch_x=-24 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C307 N$1065 N$1067 N$1111 N$1082 "Waveguide Crossing" sch_x=-22 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C308 N$1069 N$1071 N$1084 N$1086 "Waveguide Crossing" sch_x=-22 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C309 N$1073 N$1075 N$1088 N$1090 "Waveguide Crossing" sch_x=-22 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C310 N$1077 N$1079 N$1092 N$1125 "Waveguide Crossing" sch_x=-22 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C311 N$1081 N$1083 N$1113 N$1094 "Waveguide Crossing" sch_x=-20 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C312 N$1085 N$1087 N$1096 N$1098 "Waveguide Crossing" sch_x=-20 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C313 N$1089 N$1091 N$1100 N$1123 "Waveguide Crossing" sch_x=-20 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C314 N$1093 N$1095 N$1115 N$1102 "Waveguide Crossing" sch_x=-18 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C315 N$1097 N$1099 N$1104 N$1121 "Waveguide Crossing" sch_x=-18 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C316 N$1101 N$1103 N$1117 N$1119 "Waveguide Crossing" sch_x=-16 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S261 N$1120 N$1122 N$949 N$914 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S262 N$1124 N$1126 N$916 N$918 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S263 N$1128 N$1130 N$920 N$922 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S264 N$1132 N$1136 N$924 N$951 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C265 N$913 N$915 N$937 N$926 "Waveguide Crossing" sch_x=-12 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C266 N$917 N$919 N$928 N$930 "Waveguide Crossing" sch_x=-12 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C267 N$921 N$923 N$932 N$947 "Waveguide Crossing" sch_x=-12 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C268 N$925 N$927 N$939 N$934 "Waveguide Crossing" sch_x=-10 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C269 N$929 N$931 N$936 N$945 "Waveguide Crossing" sch_x=-10 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C270 N$933 N$935 N$941 N$943 "Waveguide Crossing" sch_x=-8 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S209 N$1134 N$1106 N$773 N$738 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S210 N$1108 N$1110 N$740 N$742 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S211 N$1112 N$1114 N$744 N$746 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S212 N$1116 N$1118 N$748 N$775 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C213 N$737 N$739 N$761 N$750 "Waveguide Crossing" sch_x=-12 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C214 N$741 N$743 N$752 N$754 "Waveguide Crossing" sch_x=-12 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C215 N$745 N$747 N$756 N$771 "Waveguide Crossing" sch_x=-12 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C216 N$749 N$751 N$763 N$758 "Waveguide Crossing" sch_x=-10 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C217 N$753 N$755 N$760 N$769 "Waveguide Crossing" sch_x=-10 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C218 N$757 N$759 N$765 N$767 "Waveguide Crossing" sch_x=-8 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S105 N$1822 N$1762 N$493 N$354 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S106 N$1764 N$1766 N$356 N$358 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S107 N$1768 N$1770 N$360 N$362 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S108 N$1772 N$1774 N$364 N$366 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S109 N$1776 N$1778 N$368 N$370 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S110 N$1780 N$1782 N$372 N$374 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S111 N$1784 N$1786 N$376 N$378 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S112 N$1788 N$1790 N$380 N$495 BDC_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C113 N$353 N$355 N$465 N$382 "Waveguide Crossing" sch_x=-28 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C114 N$357 N$359 N$384 N$386 "Waveguide Crossing" sch_x=-28 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C115 N$361 N$363 N$388 N$390 "Waveguide Crossing" sch_x=-28 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C116 N$365 N$367 N$392 N$394 "Waveguide Crossing" sch_x=-28 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C117 N$369 N$371 N$396 N$398 "Waveguide Crossing" sch_x=-28 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C118 N$373 N$375 N$400 N$402 "Waveguide Crossing" sch_x=-28 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C119 N$377 N$379 N$404 N$491 "Waveguide Crossing" sch_x=-28 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C120 N$381 N$383 N$467 N$406 "Waveguide Crossing" sch_x=-26 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C121 N$385 N$387 N$408 N$410 "Waveguide Crossing" sch_x=-26 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C122 N$389 N$391 N$412 N$414 "Waveguide Crossing" sch_x=-26 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C123 N$393 N$395 N$416 N$418 "Waveguide Crossing" sch_x=-26 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C124 N$397 N$399 N$420 N$422 "Waveguide Crossing" sch_x=-26 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C125 N$401 N$403 N$424 N$489 "Waveguide Crossing" sch_x=-26 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C126 N$405 N$407 N$469 N$426 "Waveguide Crossing" sch_x=-24 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C127 N$409 N$411 N$428 N$430 "Waveguide Crossing" sch_x=-24 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C128 N$413 N$415 N$432 N$434 "Waveguide Crossing" sch_x=-24 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C129 N$417 N$419 N$436 N$438 "Waveguide Crossing" sch_x=-24 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C130 N$421 N$423 N$440 N$487 "Waveguide Crossing" sch_x=-24 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C131 N$425 N$427 N$471 N$442 "Waveguide Crossing" sch_x=-22 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C132 N$429 N$431 N$444 N$446 "Waveguide Crossing" sch_x=-22 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C133 N$433 N$435 N$448 N$450 "Waveguide Crossing" sch_x=-22 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C134 N$437 N$439 N$452 N$485 "Waveguide Crossing" sch_x=-22 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C135 N$441 N$443 N$473 N$454 "Waveguide Crossing" sch_x=-20 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C136 N$445 N$447 N$456 N$458 "Waveguide Crossing" sch_x=-20 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C137 N$449 N$451 N$460 N$483 "Waveguide Crossing" sch_x=-20 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C138 N$453 N$455 N$475 N$462 "Waveguide Crossing" sch_x=-18 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C139 N$457 N$459 N$464 N$481 "Waveguide Crossing" sch_x=-18 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C140 N$461 N$463 N$477 N$479 "Waveguide Crossing" sch_x=-16 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S85 N$480 N$482 N$309 N$274 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S86 N$484 N$486 N$276 N$278 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S87 N$488 N$490 N$280 N$282 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S88 N$492 N$496 N$284 N$311 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C89 N$273 N$275 N$297 N$286 "Waveguide Crossing" sch_x=-12 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C90 N$277 N$279 N$288 N$290 "Waveguide Crossing" sch_x=-12 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C91 N$281 N$283 N$292 N$307 "Waveguide Crossing" sch_x=-12 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C92 N$285 N$287 N$299 N$294 "Waveguide Crossing" sch_x=-10 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C93 N$289 N$291 N$296 N$305 "Waveguide Crossing" sch_x=-10 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C94 N$293 N$295 N$301 N$303 "Waveguide Crossing" sch_x=-8 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S33 N$494 N$466 N$133 N$98 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S34 N$468 N$470 N$100 N$102 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S35 N$472 N$474 N$104 N$106 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S36 N$476 N$478 N$108 N$135 BDC_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C37 N$97 N$99 N$121 N$110 "Waveguide Crossing" sch_x=-12 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C38 N$101 N$103 N$112 N$114 "Waveguide Crossing" sch_x=-12 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C39 N$105 N$107 N$116 N$131 "Waveguide Crossing" sch_x=-12 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C40 N$109 N$111 N$123 N$118 "Waveguide Crossing" sch_x=-10 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C41 N$113 N$115 N$120 N$129 "Waveguide Crossing" sch_x=-10 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C42 N$117 N$119 N$125 N$127 "Waveguide Crossing" sch_x=-8 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1 N$134 N$122 N$1 N$3 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2 N$124 N$126 N$5 N$11 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3 N$2401 N$2 N$13 N$15 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4 N$8 N$2402 N$17 N$23 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S5 N$2403 N$10 N$25 N$27 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6 N$12 N$2404 N$29 N$35 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S7 N$14 N$22 N$37 N$2405 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S8 N$20 N$24 N$2406 N$39 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S9 N$26 N$34 N$41 N$2407 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S10 N$32 N$36 N$2408 N$47 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S11 N$38 N$46 N$174 N$162 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S12 N$44 N$48 N$164 N$166 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C13 N$4 N$6 N$7 N$9 "Waveguide Crossing" sch_x=-4 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C14 N$16 N$18 N$21 N$19 "Waveguide Crossing" sch_x=0 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C15 N$28 N$30 N$33 N$31 "Waveguide Crossing" sch_x=0 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C16 N$40 N$42 N$45 N$43 "Waveguide Crossing" sch_x=4 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S17 N$128 N$130 N$49 N$51 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S18 N$132 N$136 N$53 N$59 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S19 N$2409 N$50 N$61 N$63 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S20 N$56 N$2410 N$65 N$71 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S21 N$2411 N$58 N$73 N$75 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S22 N$60 N$2412 N$77 N$83 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S23 N$62 N$70 N$85 N$2413 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S24 N$68 N$72 N$2414 N$87 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S25 N$74 N$82 N$89 N$2415 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S26 N$80 N$84 N$2416 N$95 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S27 N$86 N$94 N$168 N$170 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S28 N$92 N$96 N$172 N$176 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C29 N$52 N$54 N$55 N$57 "Waveguide Crossing" sch_x=-4 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C30 N$64 N$66 N$69 N$67 "Waveguide Crossing" sch_x=0 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C31 N$76 N$78 N$81 N$79 "Waveguide Crossing" sch_x=0 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C32 N$88 N$90 N$93 N$91 "Waveguide Crossing" sch_x=4 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C47 N$161 N$150 N$137 N$139 "Waveguide Crossing" sch_x=12 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C48 N$152 N$154 N$141 N$143 "Waveguide Crossing" sch_x=12 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C49 N$156 N$171 N$145 N$147 "Waveguide Crossing" sch_x=12 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C50 N$163 N$158 N$149 N$151 "Waveguide Crossing" sch_x=10 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C51 N$160 N$169 N$153 N$155 "Waveguide Crossing" sch_x=10 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C52 N$165 N$167 N$157 N$159 "Waveguide Crossing" sch_x=8 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S43 N$173 N$138 N$638 N$610 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S44 N$140 N$142 N$612 N$614 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S45 N$144 N$146 N$616 N$618 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S46 N$148 N$175 N$620 N$622 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S53 N$310 N$298 N$177 N$179 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S54 N$300 N$302 N$181 N$187 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S55 N$2417 N$178 N$189 N$191 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S56 N$184 N$2418 N$193 N$199 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S57 N$2419 N$186 N$201 N$203 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S58 N$188 N$2420 N$205 N$211 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S59 N$190 N$198 N$213 N$2421 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S60 N$196 N$200 N$2422 N$215 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S61 N$202 N$210 N$217 N$2423 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S62 N$208 N$212 N$2424 N$223 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S63 N$214 N$222 N$350 N$338 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S64 N$220 N$224 N$340 N$342 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C65 N$180 N$182 N$183 N$185 "Waveguide Crossing" sch_x=-4 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C66 N$192 N$194 N$197 N$195 "Waveguide Crossing" sch_x=0 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C67 N$204 N$206 N$209 N$207 "Waveguide Crossing" sch_x=0 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C68 N$216 N$218 N$221 N$219 "Waveguide Crossing" sch_x=4 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S69 N$304 N$306 N$225 N$227 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S70 N$308 N$312 N$229 N$235 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S71 N$2425 N$226 N$237 N$239 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S72 N$232 N$2426 N$241 N$247 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S73 N$2427 N$234 N$249 N$251 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S74 N$236 N$2428 N$253 N$259 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S75 N$238 N$246 N$261 N$2429 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S76 N$244 N$248 N$2430 N$263 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S77 N$250 N$258 N$265 N$2431 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S78 N$256 N$260 N$2432 N$271 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S79 N$262 N$270 N$344 N$346 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S80 N$268 N$272 N$348 N$352 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C81 N$228 N$230 N$231 N$233 "Waveguide Crossing" sch_x=-4 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C82 N$240 N$242 N$245 N$243 "Waveguide Crossing" sch_x=0 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C83 N$252 N$254 N$257 N$255 "Waveguide Crossing" sch_x=0 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C84 N$264 N$266 N$269 N$267 "Waveguide Crossing" sch_x=4 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C99 N$337 N$326 N$313 N$315 "Waveguide Crossing" sch_x=12 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C100 N$328 N$330 N$317 N$319 "Waveguide Crossing" sch_x=12 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C101 N$332 N$347 N$321 N$323 "Waveguide Crossing" sch_x=12 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C102 N$339 N$334 N$325 N$327 "Waveguide Crossing" sch_x=10 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C103 N$336 N$345 N$329 N$331 "Waveguide Crossing" sch_x=10 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C104 N$341 N$343 N$333 N$335 "Waveguide Crossing" sch_x=8 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S95 N$349 N$314 N$624 N$626 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S96 N$316 N$318 N$628 N$630 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S97 N$320 N$322 N$632 N$634 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S98 N$324 N$351 N$636 N$640 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C149 N$609 N$526 N$497 N$499 "Waveguide Crossing" sch_x=28 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C150 N$528 N$530 N$501 N$503 "Waveguide Crossing" sch_x=28 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C151 N$532 N$534 N$505 N$507 "Waveguide Crossing" sch_x=28 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C152 N$536 N$538 N$509 N$511 "Waveguide Crossing" sch_x=28 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C153 N$540 N$542 N$513 N$515 "Waveguide Crossing" sch_x=28 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C154 N$544 N$546 N$517 N$519 "Waveguide Crossing" sch_x=28 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C155 N$548 N$635 N$521 N$523 "Waveguide Crossing" sch_x=28 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C156 N$611 N$550 N$525 N$527 "Waveguide Crossing" sch_x=26 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C157 N$552 N$554 N$529 N$531 "Waveguide Crossing" sch_x=26 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C158 N$556 N$558 N$533 N$535 "Waveguide Crossing" sch_x=26 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C159 N$560 N$562 N$537 N$539 "Waveguide Crossing" sch_x=26 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C160 N$564 N$566 N$541 N$543 "Waveguide Crossing" sch_x=26 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C161 N$568 N$633 N$545 N$547 "Waveguide Crossing" sch_x=26 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C162 N$613 N$570 N$549 N$551 "Waveguide Crossing" sch_x=24 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C163 N$572 N$574 N$553 N$555 "Waveguide Crossing" sch_x=24 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C164 N$576 N$578 N$557 N$559 "Waveguide Crossing" sch_x=24 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C165 N$580 N$582 N$561 N$563 "Waveguide Crossing" sch_x=24 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C166 N$584 N$631 N$565 N$567 "Waveguide Crossing" sch_x=24 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C167 N$615 N$586 N$569 N$571 "Waveguide Crossing" sch_x=22 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C168 N$588 N$590 N$573 N$575 "Waveguide Crossing" sch_x=22 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C169 N$592 N$594 N$577 N$579 "Waveguide Crossing" sch_x=22 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C170 N$596 N$629 N$581 N$583 "Waveguide Crossing" sch_x=22 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C171 N$617 N$598 N$585 N$587 "Waveguide Crossing" sch_x=20 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C172 N$600 N$602 N$589 N$591 "Waveguide Crossing" sch_x=20 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C173 N$604 N$627 N$593 N$595 "Waveguide Crossing" sch_x=20 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C174 N$619 N$606 N$597 N$599 "Waveguide Crossing" sch_x=18 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C175 N$608 N$625 N$601 N$603 "Waveguide Crossing" sch_x=18 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C176 N$621 N$623 N$605 N$607 "Waveguide Crossing" sch_x=16 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S141 N$637 N$498 N$2366 N$2306 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S142 N$500 N$502 N$2308 N$2310 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S143 N$504 N$506 N$2312 N$2314 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S144 N$508 N$510 N$2316 N$2318 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S145 N$512 N$514 N$2320 N$2322 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S146 N$516 N$518 N$2324 N$2326 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S147 N$520 N$522 N$2328 N$2330 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S148 N$524 N$639 N$2332 N$2334 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S177 N$774 N$762 N$641 N$643 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S178 N$764 N$766 N$645 N$651 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S179 N$2433 N$642 N$653 N$655 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S180 N$648 N$2434 N$657 N$663 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S181 N$2435 N$650 N$665 N$667 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S182 N$652 N$2436 N$669 N$675 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S183 N$654 N$662 N$677 N$2437 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S184 N$660 N$664 N$2438 N$679 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S185 N$666 N$674 N$681 N$2439 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S186 N$672 N$676 N$2440 N$687 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S187 N$678 N$686 N$814 N$802 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S188 N$684 N$688 N$804 N$806 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C189 N$644 N$646 N$647 N$649 "Waveguide Crossing" sch_x=-4 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C190 N$656 N$658 N$661 N$659 "Waveguide Crossing" sch_x=0 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C191 N$668 N$670 N$673 N$671 "Waveguide Crossing" sch_x=0 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C192 N$680 N$682 N$685 N$683 "Waveguide Crossing" sch_x=4 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S193 N$768 N$770 N$689 N$691 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S194 N$772 N$776 N$693 N$699 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S195 N$2441 N$690 N$701 N$703 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S196 N$696 N$2442 N$705 N$711 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S197 N$2443 N$698 N$713 N$715 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S198 N$700 N$2444 N$717 N$723 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S199 N$702 N$710 N$725 N$2445 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S200 N$708 N$712 N$2446 N$727 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S201 N$714 N$722 N$729 N$2447 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S202 N$720 N$724 N$2448 N$735 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S203 N$726 N$734 N$808 N$810 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S204 N$732 N$736 N$812 N$816 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C205 N$692 N$694 N$695 N$697 "Waveguide Crossing" sch_x=-4 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C206 N$704 N$706 N$709 N$707 "Waveguide Crossing" sch_x=0 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C207 N$716 N$718 N$721 N$719 "Waveguide Crossing" sch_x=0 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C208 N$728 N$730 N$733 N$731 "Waveguide Crossing" sch_x=4 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C223 N$801 N$790 N$777 N$779 "Waveguide Crossing" sch_x=12 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C224 N$792 N$794 N$781 N$783 "Waveguide Crossing" sch_x=12 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C225 N$796 N$811 N$785 N$787 "Waveguide Crossing" sch_x=12 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C226 N$803 N$798 N$789 N$791 "Waveguide Crossing" sch_x=10 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C227 N$800 N$809 N$793 N$795 "Waveguide Crossing" sch_x=10 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C228 N$805 N$807 N$797 N$799 "Waveguide Crossing" sch_x=8 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S219 N$813 N$778 N$1278 N$1250 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S220 N$780 N$782 N$1252 N$1254 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S221 N$784 N$786 N$1256 N$1258 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S222 N$788 N$815 N$1260 N$1262 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S229 N$950 N$938 N$817 N$819 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S230 N$940 N$942 N$821 N$827 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S231 N$2449 N$818 N$829 N$831 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S232 N$824 N$2450 N$833 N$839 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S233 N$2451 N$826 N$841 N$843 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S234 N$828 N$2452 N$845 N$851 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S235 N$830 N$838 N$853 N$2453 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S236 N$836 N$840 N$2454 N$855 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S237 N$842 N$850 N$857 N$2455 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S238 N$848 N$852 N$2456 N$863 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S239 N$854 N$862 N$990 N$978 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S240 N$860 N$864 N$980 N$982 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C241 N$820 N$822 N$823 N$825 "Waveguide Crossing" sch_x=-4 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C242 N$832 N$834 N$837 N$835 "Waveguide Crossing" sch_x=0 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C243 N$844 N$846 N$849 N$847 "Waveguide Crossing" sch_x=0 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C244 N$856 N$858 N$861 N$859 "Waveguide Crossing" sch_x=4 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S245 N$944 N$946 N$865 N$867 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S246 N$948 N$952 N$869 N$875 BDC_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S247 N$2457 N$866 N$877 N$879 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S248 N$872 N$2458 N$881 N$887 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S249 N$2459 N$874 N$889 N$891 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S250 N$876 N$2460 N$893 N$899 BDC_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S251 N$878 N$886 N$901 N$2461 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S252 N$884 N$888 N$2462 N$903 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S253 N$890 N$898 N$905 N$2463 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S254 N$896 N$900 N$2464 N$911 BDC_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S255 N$902 N$910 N$984 N$986 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S256 N$908 N$912 N$988 N$992 BDC_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C257 N$868 N$870 N$871 N$873 "Waveguide Crossing" sch_x=-4 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C258 N$880 N$882 N$885 N$883 "Waveguide Crossing" sch_x=0 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C259 N$892 N$894 N$897 N$895 "Waveguide Crossing" sch_x=0 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C260 N$904 N$906 N$909 N$907 "Waveguide Crossing" sch_x=4 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C275 N$977 N$966 N$953 N$955 "Waveguide Crossing" sch_x=12 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C276 N$968 N$970 N$957 N$959 "Waveguide Crossing" sch_x=12 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C277 N$972 N$987 N$961 N$963 "Waveguide Crossing" sch_x=12 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C278 N$979 N$974 N$965 N$967 "Waveguide Crossing" sch_x=10 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C279 N$976 N$985 N$969 N$971 "Waveguide Crossing" sch_x=10 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C280 N$981 N$983 N$973 N$975 "Waveguide Crossing" sch_x=8 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S271 N$989 N$954 N$1264 N$1266 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S272 N$956 N$958 N$1268 N$1270 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S273 N$960 N$962 N$1272 N$1274 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S274 N$964 N$991 N$1276 N$1280 BDC_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C325 N$1249 N$1166 N$1137 N$1139 "Waveguide Crossing" sch_x=28 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C326 N$1168 N$1170 N$1141 N$1143 "Waveguide Crossing" sch_x=28 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C327 N$1172 N$1174 N$1145 N$1147 "Waveguide Crossing" sch_x=28 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C328 N$1176 N$1178 N$1149 N$1151 "Waveguide Crossing" sch_x=28 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C329 N$1180 N$1182 N$1153 N$1155 "Waveguide Crossing" sch_x=28 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C330 N$1184 N$1186 N$1157 N$1159 "Waveguide Crossing" sch_x=28 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C331 N$1188 N$1275 N$1161 N$1163 "Waveguide Crossing" sch_x=28 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C332 N$1251 N$1190 N$1165 N$1167 "Waveguide Crossing" sch_x=26 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C333 N$1192 N$1194 N$1169 N$1171 "Waveguide Crossing" sch_x=26 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C334 N$1196 N$1198 N$1173 N$1175 "Waveguide Crossing" sch_x=26 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C335 N$1200 N$1202 N$1177 N$1179 "Waveguide Crossing" sch_x=26 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C336 N$1204 N$1206 N$1181 N$1183 "Waveguide Crossing" sch_x=26 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C337 N$1208 N$1273 N$1185 N$1187 "Waveguide Crossing" sch_x=26 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C338 N$1253 N$1210 N$1189 N$1191 "Waveguide Crossing" sch_x=24 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C339 N$1212 N$1214 N$1193 N$1195 "Waveguide Crossing" sch_x=24 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C340 N$1216 N$1218 N$1197 N$1199 "Waveguide Crossing" sch_x=24 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C341 N$1220 N$1222 N$1201 N$1203 "Waveguide Crossing" sch_x=24 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C342 N$1224 N$1271 N$1205 N$1207 "Waveguide Crossing" sch_x=24 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C343 N$1255 N$1226 N$1209 N$1211 "Waveguide Crossing" sch_x=22 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C344 N$1228 N$1230 N$1213 N$1215 "Waveguide Crossing" sch_x=22 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C345 N$1232 N$1234 N$1217 N$1219 "Waveguide Crossing" sch_x=22 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C346 N$1236 N$1269 N$1221 N$1223 "Waveguide Crossing" sch_x=22 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C347 N$1257 N$1238 N$1225 N$1227 "Waveguide Crossing" sch_x=20 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C348 N$1240 N$1242 N$1229 N$1231 "Waveguide Crossing" sch_x=20 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C349 N$1244 N$1267 N$1233 N$1235 "Waveguide Crossing" sch_x=20 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C350 N$1259 N$1246 N$1237 N$1239 "Waveguide Crossing" sch_x=18 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C351 N$1248 N$1265 N$1241 N$1243 "Waveguide Crossing" sch_x=18 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C352 N$1261 N$1263 N$1245 N$1247 "Waveguide Crossing" sch_x=16 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S317 N$1277 N$1138 N$2336 N$2338 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S318 N$1140 N$1142 N$2340 N$2342 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S319 N$1144 N$1146 N$2344 N$2346 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S320 N$1148 N$1150 N$2348 N$2350 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S321 N$1152 N$1154 N$2352 N$2354 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S322 N$1156 N$1158 N$2356 N$2358 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S323 N$1160 N$1162 N$2360 N$2362 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S324 N$1164 N$1279 N$2364 N$2368 BDC_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C505 N$2305 N$1886 N$1825 N$1827 "Waveguide Crossing" sch_x=60 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C506 N$1888 N$1890 N$1829 N$1831 "Waveguide Crossing" sch_x=60 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C507 N$1892 N$1894 N$1833 N$1835 "Waveguide Crossing" sch_x=60 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C508 N$1896 N$1898 N$1837 N$1839 "Waveguide Crossing" sch_x=60 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C509 N$1900 N$1902 N$1841 N$1843 "Waveguide Crossing" sch_x=60 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C510 N$1904 N$1906 N$1845 N$1847 "Waveguide Crossing" sch_x=60 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C511 N$1908 N$1910 N$1849 N$1851 "Waveguide Crossing" sch_x=60 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C512 N$1912 N$1914 N$1853 N$1855 "Waveguide Crossing" sch_x=60 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C513 N$1916 N$1918 N$1857 N$1859 "Waveguide Crossing" sch_x=60 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C514 N$1920 N$1922 N$1861 N$1863 "Waveguide Crossing" sch_x=60 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C515 N$1924 N$1926 N$1865 N$1867 "Waveguide Crossing" sch_x=60 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C516 N$1928 N$1930 N$1869 N$1871 "Waveguide Crossing" sch_x=60 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C517 N$1932 N$1934 N$1873 N$1875 "Waveguide Crossing" sch_x=60 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C518 N$1936 N$1938 N$1877 N$1879 "Waveguide Crossing" sch_x=60 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C519 N$1940 N$2363 N$1881 N$1883 "Waveguide Crossing" sch_x=60 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C520 N$2307 N$1942 N$1885 N$1887 "Waveguide Crossing" sch_x=58 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C521 N$1944 N$1946 N$1889 N$1891 "Waveguide Crossing" sch_x=58 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C522 N$1948 N$1950 N$1893 N$1895 "Waveguide Crossing" sch_x=58 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C523 N$1952 N$1954 N$1897 N$1899 "Waveguide Crossing" sch_x=58 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C524 N$1956 N$1958 N$1901 N$1903 "Waveguide Crossing" sch_x=58 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C525 N$1960 N$1962 N$1905 N$1907 "Waveguide Crossing" sch_x=58 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C526 N$1964 N$1966 N$1909 N$1911 "Waveguide Crossing" sch_x=58 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C527 N$1968 N$1970 N$1913 N$1915 "Waveguide Crossing" sch_x=58 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C528 N$1972 N$1974 N$1917 N$1919 "Waveguide Crossing" sch_x=58 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C529 N$1976 N$1978 N$1921 N$1923 "Waveguide Crossing" sch_x=58 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C530 N$1980 N$1982 N$1925 N$1927 "Waveguide Crossing" sch_x=58 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C531 N$1984 N$1986 N$1929 N$1931 "Waveguide Crossing" sch_x=58 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C532 N$1988 N$1990 N$1933 N$1935 "Waveguide Crossing" sch_x=58 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C533 N$1992 N$2361 N$1937 N$1939 "Waveguide Crossing" sch_x=58 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C534 N$2309 N$1994 N$1941 N$1943 "Waveguide Crossing" sch_x=56 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C535 N$1996 N$1998 N$1945 N$1947 "Waveguide Crossing" sch_x=56 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C536 N$2000 N$2002 N$1949 N$1951 "Waveguide Crossing" sch_x=56 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C537 N$2004 N$2006 N$1953 N$1955 "Waveguide Crossing" sch_x=56 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C538 N$2008 N$2010 N$1957 N$1959 "Waveguide Crossing" sch_x=56 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C539 N$2012 N$2014 N$1961 N$1963 "Waveguide Crossing" sch_x=56 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C540 N$2016 N$2018 N$1965 N$1967 "Waveguide Crossing" sch_x=56 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C541 N$2020 N$2022 N$1969 N$1971 "Waveguide Crossing" sch_x=56 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C542 N$2024 N$2026 N$1973 N$1975 "Waveguide Crossing" sch_x=56 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C543 N$2028 N$2030 N$1977 N$1979 "Waveguide Crossing" sch_x=56 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C544 N$2032 N$2034 N$1981 N$1983 "Waveguide Crossing" sch_x=56 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C545 N$2036 N$2038 N$1985 N$1987 "Waveguide Crossing" sch_x=56 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C546 N$2040 N$2359 N$1989 N$1991 "Waveguide Crossing" sch_x=56 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C547 N$2311 N$2042 N$1993 N$1995 "Waveguide Crossing" sch_x=54 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C548 N$2044 N$2046 N$1997 N$1999 "Waveguide Crossing" sch_x=54 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C549 N$2048 N$2050 N$2001 N$2003 "Waveguide Crossing" sch_x=54 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C550 N$2052 N$2054 N$2005 N$2007 "Waveguide Crossing" sch_x=54 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C551 N$2056 N$2058 N$2009 N$2011 "Waveguide Crossing" sch_x=54 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C552 N$2060 N$2062 N$2013 N$2015 "Waveguide Crossing" sch_x=54 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C553 N$2064 N$2066 N$2017 N$2019 "Waveguide Crossing" sch_x=54 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C554 N$2068 N$2070 N$2021 N$2023 "Waveguide Crossing" sch_x=54 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C555 N$2072 N$2074 N$2025 N$2027 "Waveguide Crossing" sch_x=54 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C556 N$2076 N$2078 N$2029 N$2031 "Waveguide Crossing" sch_x=54 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C557 N$2080 N$2082 N$2033 N$2035 "Waveguide Crossing" sch_x=54 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C558 N$2084 N$2357 N$2037 N$2039 "Waveguide Crossing" sch_x=54 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C559 N$2313 N$2086 N$2041 N$2043 "Waveguide Crossing" sch_x=52 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C560 N$2088 N$2090 N$2045 N$2047 "Waveguide Crossing" sch_x=52 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C561 N$2092 N$2094 N$2049 N$2051 "Waveguide Crossing" sch_x=52 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C562 N$2096 N$2098 N$2053 N$2055 "Waveguide Crossing" sch_x=52 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C563 N$2100 N$2102 N$2057 N$2059 "Waveguide Crossing" sch_x=52 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C564 N$2104 N$2106 N$2061 N$2063 "Waveguide Crossing" sch_x=52 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C565 N$2108 N$2110 N$2065 N$2067 "Waveguide Crossing" sch_x=52 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C566 N$2112 N$2114 N$2069 N$2071 "Waveguide Crossing" sch_x=52 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C567 N$2116 N$2118 N$2073 N$2075 "Waveguide Crossing" sch_x=52 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C568 N$2120 N$2122 N$2077 N$2079 "Waveguide Crossing" sch_x=52 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C569 N$2124 N$2355 N$2081 N$2083 "Waveguide Crossing" sch_x=52 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C570 N$2315 N$2126 N$2085 N$2087 "Waveguide Crossing" sch_x=50 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C571 N$2128 N$2130 N$2089 N$2091 "Waveguide Crossing" sch_x=50 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C572 N$2132 N$2134 N$2093 N$2095 "Waveguide Crossing" sch_x=50 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C573 N$2136 N$2138 N$2097 N$2099 "Waveguide Crossing" sch_x=50 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C574 N$2140 N$2142 N$2101 N$2103 "Waveguide Crossing" sch_x=50 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C575 N$2144 N$2146 N$2105 N$2107 "Waveguide Crossing" sch_x=50 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C576 N$2148 N$2150 N$2109 N$2111 "Waveguide Crossing" sch_x=50 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C577 N$2152 N$2154 N$2113 N$2115 "Waveguide Crossing" sch_x=50 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C578 N$2156 N$2158 N$2117 N$2119 "Waveguide Crossing" sch_x=50 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C579 N$2160 N$2353 N$2121 N$2123 "Waveguide Crossing" sch_x=50 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C580 N$2317 N$2162 N$2125 N$2127 "Waveguide Crossing" sch_x=48 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C581 N$2164 N$2166 N$2129 N$2131 "Waveguide Crossing" sch_x=48 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C582 N$2168 N$2170 N$2133 N$2135 "Waveguide Crossing" sch_x=48 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C583 N$2172 N$2174 N$2137 N$2139 "Waveguide Crossing" sch_x=48 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C584 N$2176 N$2178 N$2141 N$2143 "Waveguide Crossing" sch_x=48 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C585 N$2180 N$2182 N$2145 N$2147 "Waveguide Crossing" sch_x=48 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C586 N$2184 N$2186 N$2149 N$2151 "Waveguide Crossing" sch_x=48 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C587 N$2188 N$2190 N$2153 N$2155 "Waveguide Crossing" sch_x=48 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C588 N$2192 N$2351 N$2157 N$2159 "Waveguide Crossing" sch_x=48 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C589 N$2319 N$2194 N$2161 N$2163 "Waveguide Crossing" sch_x=46 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C590 N$2196 N$2198 N$2165 N$2167 "Waveguide Crossing" sch_x=46 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C591 N$2200 N$2202 N$2169 N$2171 "Waveguide Crossing" sch_x=46 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C592 N$2204 N$2206 N$2173 N$2175 "Waveguide Crossing" sch_x=46 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C593 N$2208 N$2210 N$2177 N$2179 "Waveguide Crossing" sch_x=46 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C594 N$2212 N$2214 N$2181 N$2183 "Waveguide Crossing" sch_x=46 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C595 N$2216 N$2218 N$2185 N$2187 "Waveguide Crossing" sch_x=46 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C596 N$2220 N$2349 N$2189 N$2191 "Waveguide Crossing" sch_x=46 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C597 N$2321 N$2222 N$2193 N$2195 "Waveguide Crossing" sch_x=44 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C598 N$2224 N$2226 N$2197 N$2199 "Waveguide Crossing" sch_x=44 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C599 N$2228 N$2230 N$2201 N$2203 "Waveguide Crossing" sch_x=44 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C600 N$2232 N$2234 N$2205 N$2207 "Waveguide Crossing" sch_x=44 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C601 N$2236 N$2238 N$2209 N$2211 "Waveguide Crossing" sch_x=44 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C602 N$2240 N$2242 N$2213 N$2215 "Waveguide Crossing" sch_x=44 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C603 N$2244 N$2347 N$2217 N$2219 "Waveguide Crossing" sch_x=44 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C604 N$2323 N$2246 N$2221 N$2223 "Waveguide Crossing" sch_x=42 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C605 N$2248 N$2250 N$2225 N$2227 "Waveguide Crossing" sch_x=42 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C606 N$2252 N$2254 N$2229 N$2231 "Waveguide Crossing" sch_x=42 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C607 N$2256 N$2258 N$2233 N$2235 "Waveguide Crossing" sch_x=42 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C608 N$2260 N$2262 N$2237 N$2239 "Waveguide Crossing" sch_x=42 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C609 N$2264 N$2345 N$2241 N$2243 "Waveguide Crossing" sch_x=42 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C610 N$2325 N$2266 N$2245 N$2247 "Waveguide Crossing" sch_x=40 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C611 N$2268 N$2270 N$2249 N$2251 "Waveguide Crossing" sch_x=40 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C612 N$2272 N$2274 N$2253 N$2255 "Waveguide Crossing" sch_x=40 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C613 N$2276 N$2278 N$2257 N$2259 "Waveguide Crossing" sch_x=40 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C614 N$2280 N$2343 N$2261 N$2263 "Waveguide Crossing" sch_x=40 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C615 N$2327 N$2282 N$2265 N$2267 "Waveguide Crossing" sch_x=38 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C616 N$2284 N$2286 N$2269 N$2271 "Waveguide Crossing" sch_x=38 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C617 N$2288 N$2290 N$2273 N$2275 "Waveguide Crossing" sch_x=38 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C618 N$2292 N$2341 N$2277 N$2279 "Waveguide Crossing" sch_x=38 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C619 N$2329 N$2294 N$2281 N$2283 "Waveguide Crossing" sch_x=36 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C620 N$2296 N$2298 N$2285 N$2287 "Waveguide Crossing" sch_x=36 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C621 N$2300 N$2339 N$2289 N$2291 "Waveguide Crossing" sch_x=36 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C622 N$2331 N$2302 N$2293 N$2295 "Waveguide Crossing" sch_x=34 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C623 N$2304 N$2337 N$2297 N$2299 "Waveguide Crossing" sch_x=34 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C624 N$2333 N$2335 N$2301 N$2303 "Waveguide Crossing" sch_x=32 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S489 N$2365 N$1826 N$2465 N$2466 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S490 N$1828 N$1830 N$2467 N$2468 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S491 N$1832 N$1834 N$2469 N$2470 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S492 N$1836 N$1838 N$2471 N$2472 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S493 N$1840 N$1842 N$2473 N$2474 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S494 N$1844 N$1846 N$2475 N$2476 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S495 N$1848 N$1850 N$2477 N$2478 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S496 N$1852 N$1854 N$2479 N$2480 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S497 N$1856 N$1858 N$2481 N$2482 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S498 N$1860 N$1862 N$2483 N$2484 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S499 N$1864 N$1866 N$2485 N$2486 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S500 N$1868 N$1870 N$2487 N$2488 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S501 N$1872 N$1874 N$2489 N$2490 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S502 N$1876 N$1878 N$2491 N$2492 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S503 N$1880 N$1882 N$2493 N$2494 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S504 N$1884 N$2367 N$2495 N$2496 BDC_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1 N$1 N$2 "Straight Waveguide" sch_x=-4 sch_y=15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2 N$3 N$4 "Straight Waveguide" sch_x=-5 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3 N$5 N$6 "Straight Waveguide" sch_x=-5 sch_y=13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4 N$7 N$8 "Straight Waveguide" sch_x=-3 sch_y=14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5 N$9 N$10 "Straight Waveguide" sch_x=-3 sch_y=13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6 N$11 N$12 "Straight Waveguide" sch_x=-4 sch_y=12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7 N$13 N$14 "Straight Waveguide" sch_x=0 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8 N$15 N$16 "Straight Waveguide" sch_x=-1 sch_y=15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9 N$17 N$18 "Straight Waveguide" sch_x=-1 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10 N$19 N$20 "Straight Waveguide" sch_x=1 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11 N$21 N$22 "Straight Waveguide" sch_x=1 sch_y=15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12 N$23 N$24 "Straight Waveguide" sch_x=0 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13 N$25 N$26 "Straight Waveguide" sch_x=0 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14 N$27 N$28 "Straight Waveguide" sch_x=-1 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15 N$29 N$30 "Straight Waveguide" sch_x=-1 sch_y=12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16 N$31 N$32 "Straight Waveguide" sch_x=1 sch_y=12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17 N$33 N$34 "Straight Waveguide" sch_x=1 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W18 N$35 N$36 "Straight Waveguide" sch_x=0 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W19 N$37 N$38 "Straight Waveguide" sch_x=4 sch_y=15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W20 N$39 N$40 "Straight Waveguide" sch_x=3 sch_y=14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W21 N$41 N$42 "Straight Waveguide" sch_x=3 sch_y=13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W22 N$43 N$44 "Straight Waveguide" sch_x=5 sch_y=13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W23 N$45 N$46 "Straight Waveguide" sch_x=5 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W24 N$47 N$48 "Straight Waveguide" sch_x=4 sch_y=12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W25 N$49 N$50 "Straight Waveguide" sch_x=-4 sch_y=11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W26 N$51 N$52 "Straight Waveguide" sch_x=-5 sch_y=10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W27 N$53 N$54 "Straight Waveguide" sch_x=-5 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W28 N$55 N$56 "Straight Waveguide" sch_x=-3 sch_y=10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W29 N$57 N$58 "Straight Waveguide" sch_x=-3 sch_y=9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W30 N$59 N$60 "Straight Waveguide" sch_x=-4 sch_y=8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W31 N$61 N$62 "Straight Waveguide" sch_x=0 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W32 N$63 N$64 "Straight Waveguide" sch_x=-1 sch_y=11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W33 N$65 N$66 "Straight Waveguide" sch_x=-1 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W34 N$67 N$68 "Straight Waveguide" sch_x=1 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W35 N$69 N$70 "Straight Waveguide" sch_x=1 sch_y=11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W36 N$71 N$72 "Straight Waveguide" sch_x=0 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W37 N$73 N$74 "Straight Waveguide" sch_x=0 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W38 N$75 N$76 "Straight Waveguide" sch_x=-1 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W39 N$77 N$78 "Straight Waveguide" sch_x=-1 sch_y=8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W40 N$79 N$80 "Straight Waveguide" sch_x=1 sch_y=8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W41 N$81 N$82 "Straight Waveguide" sch_x=1 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W42 N$83 N$84 "Straight Waveguide" sch_x=0 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W43 N$85 N$86 "Straight Waveguide" sch_x=4 sch_y=11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W44 N$87 N$88 "Straight Waveguide" sch_x=3 sch_y=10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W45 N$89 N$90 "Straight Waveguide" sch_x=3 sch_y=9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W46 N$91 N$92 "Straight Waveguide" sch_x=5 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W47 N$93 N$94 "Straight Waveguide" sch_x=5 sch_y=10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W48 N$95 N$96 "Straight Waveguide" sch_x=4 sch_y=8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W49 N$98 N$97 "Straight Waveguide" sch_x=-13 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W50 N$100 N$99 "Straight Waveguide" sch_x=-13 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W51 N$102 N$101 "Straight Waveguide" sch_x=-13 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W52 N$104 N$103 "Straight Waveguide" sch_x=-13 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W53 N$106 N$105 "Straight Waveguide" sch_x=-13 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W54 N$108 N$107 "Straight Waveguide" sch_x=-13 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W55 N$110 N$109 "Straight Waveguide" sch_x=-11 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W56 N$112 N$111 "Straight Waveguide" sch_x=-11 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W57 N$114 N$113 "Straight Waveguide" sch_x=-11 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W58 N$116 N$115 "Straight Waveguide" sch_x=-11 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W59 N$118 N$117 "Straight Waveguide" sch_x=-9 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W60 N$120 N$119 "Straight Waveguide" sch_x=-9 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W61 N$121 N$122 "Straight Waveguide" sch_x=-9 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W62 N$123 N$124 "Straight Waveguide" sch_x=-8 sch_y=13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W63 N$125 N$126 "Straight Waveguide" sch_x=-7 sch_y=12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W64 N$127 N$128 "Straight Waveguide" sch_x=-7 sch_y=11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W65 N$129 N$130 "Straight Waveguide" sch_x=-8 sch_y=10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W66 N$131 N$132 "Straight Waveguide" sch_x=-9 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W67 N$133 N$134 "Straight Waveguide" sch_x=-10 sch_y=14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W68 N$135 N$136 "Straight Waveguide" sch_x=-10 sch_y=9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W69 N$137 N$138 "Straight Waveguide" sch_x=13 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W70 N$139 N$140 "Straight Waveguide" sch_x=13 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W71 N$141 N$142 "Straight Waveguide" sch_x=13 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W72 N$143 N$144 "Straight Waveguide" sch_x=13 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W73 N$145 N$146 "Straight Waveguide" sch_x=13 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W74 N$147 N$148 "Straight Waveguide" sch_x=13 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W75 N$149 N$150 "Straight Waveguide" sch_x=11 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W76 N$151 N$152 "Straight Waveguide" sch_x=11 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W77 N$153 N$154 "Straight Waveguide" sch_x=11 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W78 N$155 N$156 "Straight Waveguide" sch_x=11 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W79 N$157 N$158 "Straight Waveguide" sch_x=9 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W80 N$159 N$160 "Straight Waveguide" sch_x=9 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W81 N$162 N$161 "Straight Waveguide" sch_x=9 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W82 N$164 N$163 "Straight Waveguide" sch_x=8 sch_y=13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W83 N$166 N$165 "Straight Waveguide" sch_x=7 sch_y=12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W84 N$168 N$167 "Straight Waveguide" sch_x=7 sch_y=11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W85 N$170 N$169 "Straight Waveguide" sch_x=8 sch_y=10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W86 N$172 N$171 "Straight Waveguide" sch_x=9 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W87 N$174 N$173 "Straight Waveguide" sch_x=10 sch_y=14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W88 N$176 N$175 "Straight Waveguide" sch_x=10 sch_y=9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W89 N$177 N$178 "Straight Waveguide" sch_x=-4 sch_y=7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W90 N$179 N$180 "Straight Waveguide" sch_x=-5 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W91 N$181 N$182 "Straight Waveguide" sch_x=-5 sch_y=5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W92 N$183 N$184 "Straight Waveguide" sch_x=-3 sch_y=6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W93 N$185 N$186 "Straight Waveguide" sch_x=-3 sch_y=5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W94 N$187 N$188 "Straight Waveguide" sch_x=-4 sch_y=4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W95 N$189 N$190 "Straight Waveguide" sch_x=0 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W96 N$191 N$192 "Straight Waveguide" sch_x=-1 sch_y=7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W97 N$193 N$194 "Straight Waveguide" sch_x=-1 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W98 N$195 N$196 "Straight Waveguide" sch_x=1 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W99 N$197 N$198 "Straight Waveguide" sch_x=1 sch_y=7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W100 N$199 N$200 "Straight Waveguide" sch_x=0 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W101 N$201 N$202 "Straight Waveguide" sch_x=0 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W102 N$203 N$204 "Straight Waveguide" sch_x=-1 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W103 N$205 N$206 "Straight Waveguide" sch_x=-1 sch_y=4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W104 N$207 N$208 "Straight Waveguide" sch_x=1 sch_y=4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W105 N$209 N$210 "Straight Waveguide" sch_x=1 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W106 N$211 N$212 "Straight Waveguide" sch_x=0 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W107 N$213 N$214 "Straight Waveguide" sch_x=4 sch_y=7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W108 N$215 N$216 "Straight Waveguide" sch_x=3 sch_y=6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W109 N$217 N$218 "Straight Waveguide" sch_x=3 sch_y=5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W110 N$219 N$220 "Straight Waveguide" sch_x=5 sch_y=5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W111 N$221 N$222 "Straight Waveguide" sch_x=5 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W112 N$223 N$224 "Straight Waveguide" sch_x=4 sch_y=4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W113 N$225 N$226 "Straight Waveguide" sch_x=-4 sch_y=3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W114 N$227 N$228 "Straight Waveguide" sch_x=-5 sch_y=2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W115 N$229 N$230 "Straight Waveguide" sch_x=-5 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W116 N$231 N$232 "Straight Waveguide" sch_x=-3 sch_y=2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W117 N$233 N$234 "Straight Waveguide" sch_x=-3 sch_y=1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W118 N$235 N$236 "Straight Waveguide" sch_x=-4 sch_y=0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W119 N$237 N$238 "Straight Waveguide" sch_x=0 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W120 N$239 N$240 "Straight Waveguide" sch_x=-1 sch_y=3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W121 N$241 N$242 "Straight Waveguide" sch_x=-1 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W122 N$243 N$244 "Straight Waveguide" sch_x=1 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W123 N$245 N$246 "Straight Waveguide" sch_x=1 sch_y=3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W124 N$247 N$248 "Straight Waveguide" sch_x=0 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W125 N$249 N$250 "Straight Waveguide" sch_x=0 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W126 N$251 N$252 "Straight Waveguide" sch_x=-1 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W127 N$253 N$254 "Straight Waveguide" sch_x=-1 sch_y=0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W128 N$255 N$256 "Straight Waveguide" sch_x=1 sch_y=0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W129 N$257 N$258 "Straight Waveguide" sch_x=1 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W130 N$259 N$260 "Straight Waveguide" sch_x=0 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W131 N$261 N$262 "Straight Waveguide" sch_x=4 sch_y=3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W132 N$263 N$264 "Straight Waveguide" sch_x=3 sch_y=2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W133 N$265 N$266 "Straight Waveguide" sch_x=3 sch_y=1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W134 N$267 N$268 "Straight Waveguide" sch_x=5 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W135 N$269 N$270 "Straight Waveguide" sch_x=5 sch_y=2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W136 N$271 N$272 "Straight Waveguide" sch_x=4 sch_y=0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W137 N$274 N$273 "Straight Waveguide" sch_x=-13 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W138 N$276 N$275 "Straight Waveguide" sch_x=-13 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W139 N$278 N$277 "Straight Waveguide" sch_x=-13 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W140 N$280 N$279 "Straight Waveguide" sch_x=-13 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W141 N$282 N$281 "Straight Waveguide" sch_x=-13 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W142 N$284 N$283 "Straight Waveguide" sch_x=-13 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W143 N$286 N$285 "Straight Waveguide" sch_x=-11 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W144 N$288 N$287 "Straight Waveguide" sch_x=-11 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W145 N$290 N$289 "Straight Waveguide" sch_x=-11 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W146 N$292 N$291 "Straight Waveguide" sch_x=-11 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W147 N$294 N$293 "Straight Waveguide" sch_x=-9 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W148 N$296 N$295 "Straight Waveguide" sch_x=-9 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W149 N$297 N$298 "Straight Waveguide" sch_x=-9 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W150 N$299 N$300 "Straight Waveguide" sch_x=-8 sch_y=5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W151 N$301 N$302 "Straight Waveguide" sch_x=-7 sch_y=4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W152 N$303 N$304 "Straight Waveguide" sch_x=-7 sch_y=3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W153 N$305 N$306 "Straight Waveguide" sch_x=-8 sch_y=2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W154 N$307 N$308 "Straight Waveguide" sch_x=-9 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W155 N$309 N$310 "Straight Waveguide" sch_x=-10 sch_y=6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W156 N$311 N$312 "Straight Waveguide" sch_x=-10 sch_y=1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W157 N$313 N$314 "Straight Waveguide" sch_x=13 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W158 N$315 N$316 "Straight Waveguide" sch_x=13 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W159 N$317 N$318 "Straight Waveguide" sch_x=13 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W160 N$319 N$320 "Straight Waveguide" sch_x=13 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W161 N$321 N$322 "Straight Waveguide" sch_x=13 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W162 N$323 N$324 "Straight Waveguide" sch_x=13 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W163 N$325 N$326 "Straight Waveguide" sch_x=11 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W164 N$327 N$328 "Straight Waveguide" sch_x=11 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W165 N$329 N$330 "Straight Waveguide" sch_x=11 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W166 N$331 N$332 "Straight Waveguide" sch_x=11 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W167 N$333 N$334 "Straight Waveguide" sch_x=9 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W168 N$335 N$336 "Straight Waveguide" sch_x=9 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W169 N$338 N$337 "Straight Waveguide" sch_x=9 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W170 N$340 N$339 "Straight Waveguide" sch_x=8 sch_y=5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W171 N$342 N$341 "Straight Waveguide" sch_x=7 sch_y=4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W172 N$344 N$343 "Straight Waveguide" sch_x=7 sch_y=3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W173 N$346 N$345 "Straight Waveguide" sch_x=8 sch_y=2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W174 N$348 N$347 "Straight Waveguide" sch_x=9 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W175 N$350 N$349 "Straight Waveguide" sch_x=10 sch_y=6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W176 N$352 N$351 "Straight Waveguide" sch_x=10 sch_y=1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W177 N$354 N$353 "Straight Waveguide" sch_x=-29 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W178 N$356 N$355 "Straight Waveguide" sch_x=-29 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W179 N$358 N$357 "Straight Waveguide" sch_x=-29 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W180 N$360 N$359 "Straight Waveguide" sch_x=-29 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W181 N$362 N$361 "Straight Waveguide" sch_x=-29 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W182 N$364 N$363 "Straight Waveguide" sch_x=-29 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W183 N$366 N$365 "Straight Waveguide" sch_x=-29 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W184 N$368 N$367 "Straight Waveguide" sch_x=-29 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W185 N$370 N$369 "Straight Waveguide" sch_x=-29 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W186 N$372 N$371 "Straight Waveguide" sch_x=-29 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W187 N$374 N$373 "Straight Waveguide" sch_x=-29 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W188 N$376 N$375 "Straight Waveguide" sch_x=-29 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W189 N$378 N$377 "Straight Waveguide" sch_x=-29 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W190 N$380 N$379 "Straight Waveguide" sch_x=-29 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W191 N$382 N$381 "Straight Waveguide" sch_x=-27 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W192 N$384 N$383 "Straight Waveguide" sch_x=-27 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W193 N$386 N$385 "Straight Waveguide" sch_x=-27 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W194 N$388 N$387 "Straight Waveguide" sch_x=-27 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W195 N$390 N$389 "Straight Waveguide" sch_x=-27 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W196 N$392 N$391 "Straight Waveguide" sch_x=-27 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W197 N$394 N$393 "Straight Waveguide" sch_x=-27 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W198 N$396 N$395 "Straight Waveguide" sch_x=-27 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W199 N$398 N$397 "Straight Waveguide" sch_x=-27 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W200 N$400 N$399 "Straight Waveguide" sch_x=-27 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W201 N$402 N$401 "Straight Waveguide" sch_x=-27 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W202 N$404 N$403 "Straight Waveguide" sch_x=-27 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W203 N$406 N$405 "Straight Waveguide" sch_x=-25 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W204 N$408 N$407 "Straight Waveguide" sch_x=-25 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W205 N$410 N$409 "Straight Waveguide" sch_x=-25 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W206 N$412 N$411 "Straight Waveguide" sch_x=-25 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W207 N$414 N$413 "Straight Waveguide" sch_x=-25 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W208 N$416 N$415 "Straight Waveguide" sch_x=-25 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W209 N$418 N$417 "Straight Waveguide" sch_x=-25 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W210 N$420 N$419 "Straight Waveguide" sch_x=-25 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W211 N$422 N$421 "Straight Waveguide" sch_x=-25 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W212 N$424 N$423 "Straight Waveguide" sch_x=-25 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W213 N$426 N$425 "Straight Waveguide" sch_x=-23 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W214 N$428 N$427 "Straight Waveguide" sch_x=-23 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W215 N$430 N$429 "Straight Waveguide" sch_x=-23 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W216 N$432 N$431 "Straight Waveguide" sch_x=-23 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W217 N$434 N$433 "Straight Waveguide" sch_x=-23 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W218 N$436 N$435 "Straight Waveguide" sch_x=-23 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W219 N$438 N$437 "Straight Waveguide" sch_x=-23 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W220 N$440 N$439 "Straight Waveguide" sch_x=-23 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W221 N$442 N$441 "Straight Waveguide" sch_x=-21 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W222 N$444 N$443 "Straight Waveguide" sch_x=-21 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W223 N$446 N$445 "Straight Waveguide" sch_x=-21 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W224 N$448 N$447 "Straight Waveguide" sch_x=-21 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W225 N$450 N$449 "Straight Waveguide" sch_x=-21 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W226 N$452 N$451 "Straight Waveguide" sch_x=-21 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W227 N$454 N$453 "Straight Waveguide" sch_x=-19 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W228 N$456 N$455 "Straight Waveguide" sch_x=-19 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W229 N$458 N$457 "Straight Waveguide" sch_x=-19 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W230 N$460 N$459 "Straight Waveguide" sch_x=-19 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W231 N$462 N$461 "Straight Waveguide" sch_x=-17 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W232 N$464 N$463 "Straight Waveguide" sch_x=-17 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W233 N$465 N$466 "Straight Waveguide" sch_x=-21 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W234 N$467 N$468 "Straight Waveguide" sch_x=-20 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W235 N$469 N$470 "Straight Waveguide" sch_x=-19 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W236 N$471 N$472 "Straight Waveguide" sch_x=-18 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W237 N$473 N$474 "Straight Waveguide" sch_x=-17 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W238 N$475 N$476 "Straight Waveguide" sch_x=-16 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W239 N$477 N$478 "Straight Waveguide" sch_x=-15 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W240 N$479 N$480 "Straight Waveguide" sch_x=-15 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W241 N$481 N$482 "Straight Waveguide" sch_x=-16 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W242 N$483 N$484 "Straight Waveguide" sch_x=-17 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W243 N$485 N$486 "Straight Waveguide" sch_x=-18 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W244 N$487 N$488 "Straight Waveguide" sch_x=-19 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W245 N$489 N$490 "Straight Waveguide" sch_x=-20 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W246 N$491 N$492 "Straight Waveguide" sch_x=-21 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W247 N$493 N$494 "Straight Waveguide" sch_x=-22 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W248 N$495 N$496 "Straight Waveguide" sch_x=-22 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W249 N$497 N$498 "Straight Waveguide" sch_x=29 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W250 N$499 N$500 "Straight Waveguide" sch_x=29 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W251 N$501 N$502 "Straight Waveguide" sch_x=29 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W252 N$503 N$504 "Straight Waveguide" sch_x=29 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W253 N$505 N$506 "Straight Waveguide" sch_x=29 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W254 N$507 N$508 "Straight Waveguide" sch_x=29 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W255 N$509 N$510 "Straight Waveguide" sch_x=29 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W256 N$511 N$512 "Straight Waveguide" sch_x=29 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W257 N$513 N$514 "Straight Waveguide" sch_x=29 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W258 N$515 N$516 "Straight Waveguide" sch_x=29 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W259 N$517 N$518 "Straight Waveguide" sch_x=29 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W260 N$519 N$520 "Straight Waveguide" sch_x=29 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W261 N$521 N$522 "Straight Waveguide" sch_x=29 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W262 N$523 N$524 "Straight Waveguide" sch_x=29 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W263 N$525 N$526 "Straight Waveguide" sch_x=27 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W264 N$527 N$528 "Straight Waveguide" sch_x=27 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W265 N$529 N$530 "Straight Waveguide" sch_x=27 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W266 N$531 N$532 "Straight Waveguide" sch_x=27 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W267 N$533 N$534 "Straight Waveguide" sch_x=27 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W268 N$535 N$536 "Straight Waveguide" sch_x=27 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W269 N$537 N$538 "Straight Waveguide" sch_x=27 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W270 N$539 N$540 "Straight Waveguide" sch_x=27 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W271 N$541 N$542 "Straight Waveguide" sch_x=27 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W272 N$543 N$544 "Straight Waveguide" sch_x=27 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W273 N$545 N$546 "Straight Waveguide" sch_x=27 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W274 N$547 N$548 "Straight Waveguide" sch_x=27 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W275 N$549 N$550 "Straight Waveguide" sch_x=25 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W276 N$551 N$552 "Straight Waveguide" sch_x=25 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W277 N$553 N$554 "Straight Waveguide" sch_x=25 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W278 N$555 N$556 "Straight Waveguide" sch_x=25 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W279 N$557 N$558 "Straight Waveguide" sch_x=25 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W280 N$559 N$560 "Straight Waveguide" sch_x=25 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W281 N$561 N$562 "Straight Waveguide" sch_x=25 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W282 N$563 N$564 "Straight Waveguide" sch_x=25 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W283 N$565 N$566 "Straight Waveguide" sch_x=25 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W284 N$567 N$568 "Straight Waveguide" sch_x=25 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W285 N$569 N$570 "Straight Waveguide" sch_x=23 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W286 N$571 N$572 "Straight Waveguide" sch_x=23 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W287 N$573 N$574 "Straight Waveguide" sch_x=23 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W288 N$575 N$576 "Straight Waveguide" sch_x=23 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W289 N$577 N$578 "Straight Waveguide" sch_x=23 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W290 N$579 N$580 "Straight Waveguide" sch_x=23 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W291 N$581 N$582 "Straight Waveguide" sch_x=23 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W292 N$583 N$584 "Straight Waveguide" sch_x=23 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W293 N$585 N$586 "Straight Waveguide" sch_x=21 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W294 N$587 N$588 "Straight Waveguide" sch_x=21 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W295 N$589 N$590 "Straight Waveguide" sch_x=21 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W296 N$591 N$592 "Straight Waveguide" sch_x=21 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W297 N$593 N$594 "Straight Waveguide" sch_x=21 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W298 N$595 N$596 "Straight Waveguide" sch_x=21 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W299 N$597 N$598 "Straight Waveguide" sch_x=19 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W300 N$599 N$600 "Straight Waveguide" sch_x=19 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W301 N$601 N$602 "Straight Waveguide" sch_x=19 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W302 N$603 N$604 "Straight Waveguide" sch_x=19 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W303 N$605 N$606 "Straight Waveguide" sch_x=17 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W304 N$607 N$608 "Straight Waveguide" sch_x=17 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W305 N$610 N$609 "Straight Waveguide" sch_x=21 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W306 N$612 N$611 "Straight Waveguide" sch_x=20 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W307 N$614 N$613 "Straight Waveguide" sch_x=19 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W308 N$616 N$615 "Straight Waveguide" sch_x=18 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W309 N$618 N$617 "Straight Waveguide" sch_x=17 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W310 N$620 N$619 "Straight Waveguide" sch_x=16 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W311 N$622 N$621 "Straight Waveguide" sch_x=15 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W312 N$624 N$623 "Straight Waveguide" sch_x=15 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W313 N$626 N$625 "Straight Waveguide" sch_x=16 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W314 N$628 N$627 "Straight Waveguide" sch_x=17 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W315 N$630 N$629 "Straight Waveguide" sch_x=18 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W316 N$632 N$631 "Straight Waveguide" sch_x=19 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W317 N$634 N$633 "Straight Waveguide" sch_x=20 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W318 N$636 N$635 "Straight Waveguide" sch_x=21 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W319 N$638 N$637 "Straight Waveguide" sch_x=22 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W320 N$640 N$639 "Straight Waveguide" sch_x=22 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W321 N$641 N$642 "Straight Waveguide" sch_x=-4 sch_y=-0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W322 N$643 N$644 "Straight Waveguide" sch_x=-5 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W323 N$645 N$646 "Straight Waveguide" sch_x=-5 sch_y=-2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W324 N$647 N$648 "Straight Waveguide" sch_x=-3 sch_y=-1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W325 N$649 N$650 "Straight Waveguide" sch_x=-3 sch_y=-2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W326 N$651 N$652 "Straight Waveguide" sch_x=-4 sch_y=-3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W327 N$653 N$654 "Straight Waveguide" sch_x=0 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W328 N$655 N$656 "Straight Waveguide" sch_x=-1 sch_y=-0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W329 N$657 N$658 "Straight Waveguide" sch_x=-1 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W330 N$659 N$660 "Straight Waveguide" sch_x=1 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W331 N$661 N$662 "Straight Waveguide" sch_x=1 sch_y=-0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W332 N$663 N$664 "Straight Waveguide" sch_x=0 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W333 N$665 N$666 "Straight Waveguide" sch_x=0 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W334 N$667 N$668 "Straight Waveguide" sch_x=-1 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W335 N$669 N$670 "Straight Waveguide" sch_x=-1 sch_y=-3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W336 N$671 N$672 "Straight Waveguide" sch_x=1 sch_y=-3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W337 N$673 N$674 "Straight Waveguide" sch_x=1 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W338 N$675 N$676 "Straight Waveguide" sch_x=0 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W339 N$677 N$678 "Straight Waveguide" sch_x=4 sch_y=-0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W340 N$679 N$680 "Straight Waveguide" sch_x=3 sch_y=-1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W341 N$681 N$682 "Straight Waveguide" sch_x=3 sch_y=-2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W342 N$683 N$684 "Straight Waveguide" sch_x=5 sch_y=-2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W343 N$685 N$686 "Straight Waveguide" sch_x=5 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W344 N$687 N$688 "Straight Waveguide" sch_x=4 sch_y=-3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W345 N$689 N$690 "Straight Waveguide" sch_x=-4 sch_y=-4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W346 N$691 N$692 "Straight Waveguide" sch_x=-5 sch_y=-5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W347 N$693 N$694 "Straight Waveguide" sch_x=-5 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W348 N$695 N$696 "Straight Waveguide" sch_x=-3 sch_y=-5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W349 N$697 N$698 "Straight Waveguide" sch_x=-3 sch_y=-6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W350 N$699 N$700 "Straight Waveguide" sch_x=-4 sch_y=-7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W351 N$701 N$702 "Straight Waveguide" sch_x=0 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W352 N$703 N$704 "Straight Waveguide" sch_x=-1 sch_y=-4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W353 N$705 N$706 "Straight Waveguide" sch_x=-1 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W354 N$707 N$708 "Straight Waveguide" sch_x=1 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W355 N$709 N$710 "Straight Waveguide" sch_x=1 sch_y=-4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W356 N$711 N$712 "Straight Waveguide" sch_x=0 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W357 N$713 N$714 "Straight Waveguide" sch_x=0 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W358 N$715 N$716 "Straight Waveguide" sch_x=-1 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W359 N$717 N$718 "Straight Waveguide" sch_x=-1 sch_y=-7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W360 N$719 N$720 "Straight Waveguide" sch_x=1 sch_y=-7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W361 N$721 N$722 "Straight Waveguide" sch_x=1 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W362 N$723 N$724 "Straight Waveguide" sch_x=0 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W363 N$725 N$726 "Straight Waveguide" sch_x=4 sch_y=-4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W364 N$727 N$728 "Straight Waveguide" sch_x=3 sch_y=-5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W365 N$729 N$730 "Straight Waveguide" sch_x=3 sch_y=-6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W366 N$731 N$732 "Straight Waveguide" sch_x=5 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W367 N$733 N$734 "Straight Waveguide" sch_x=5 sch_y=-5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W368 N$735 N$736 "Straight Waveguide" sch_x=4 sch_y=-7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W369 N$738 N$737 "Straight Waveguide" sch_x=-13 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W370 N$740 N$739 "Straight Waveguide" sch_x=-13 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W371 N$742 N$741 "Straight Waveguide" sch_x=-13 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W372 N$744 N$743 "Straight Waveguide" sch_x=-13 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W373 N$746 N$745 "Straight Waveguide" sch_x=-13 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W374 N$748 N$747 "Straight Waveguide" sch_x=-13 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W375 N$750 N$749 "Straight Waveguide" sch_x=-11 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W376 N$752 N$751 "Straight Waveguide" sch_x=-11 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W377 N$754 N$753 "Straight Waveguide" sch_x=-11 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W378 N$756 N$755 "Straight Waveguide" sch_x=-11 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W379 N$758 N$757 "Straight Waveguide" sch_x=-9 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W380 N$760 N$759 "Straight Waveguide" sch_x=-9 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W381 N$761 N$762 "Straight Waveguide" sch_x=-9 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W382 N$763 N$764 "Straight Waveguide" sch_x=-8 sch_y=-2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W383 N$765 N$766 "Straight Waveguide" sch_x=-7 sch_y=-3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W384 N$767 N$768 "Straight Waveguide" sch_x=-7 sch_y=-4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W385 N$769 N$770 "Straight Waveguide" sch_x=-8 sch_y=-5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W386 N$771 N$772 "Straight Waveguide" sch_x=-9 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W387 N$773 N$774 "Straight Waveguide" sch_x=-10 sch_y=-1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W388 N$775 N$776 "Straight Waveguide" sch_x=-10 sch_y=-6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W389 N$777 N$778 "Straight Waveguide" sch_x=13 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W390 N$779 N$780 "Straight Waveguide" sch_x=13 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W391 N$781 N$782 "Straight Waveguide" sch_x=13 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W392 N$783 N$784 "Straight Waveguide" sch_x=13 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W393 N$785 N$786 "Straight Waveguide" sch_x=13 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W394 N$787 N$788 "Straight Waveguide" sch_x=13 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W395 N$789 N$790 "Straight Waveguide" sch_x=11 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W396 N$791 N$792 "Straight Waveguide" sch_x=11 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W397 N$793 N$794 "Straight Waveguide" sch_x=11 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W398 N$795 N$796 "Straight Waveguide" sch_x=11 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W399 N$797 N$798 "Straight Waveguide" sch_x=9 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W400 N$799 N$800 "Straight Waveguide" sch_x=9 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W401 N$802 N$801 "Straight Waveguide" sch_x=9 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W402 N$804 N$803 "Straight Waveguide" sch_x=8 sch_y=-2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W403 N$806 N$805 "Straight Waveguide" sch_x=7 sch_y=-3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W404 N$808 N$807 "Straight Waveguide" sch_x=7 sch_y=-4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W405 N$810 N$809 "Straight Waveguide" sch_x=8 sch_y=-5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W406 N$812 N$811 "Straight Waveguide" sch_x=9 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W407 N$814 N$813 "Straight Waveguide" sch_x=10 sch_y=-1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W408 N$816 N$815 "Straight Waveguide" sch_x=10 sch_y=-6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W409 N$817 N$818 "Straight Waveguide" sch_x=-4 sch_y=-8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W410 N$819 N$820 "Straight Waveguide" sch_x=-5 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W411 N$821 N$822 "Straight Waveguide" sch_x=-5 sch_y=-10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W412 N$823 N$824 "Straight Waveguide" sch_x=-3 sch_y=-9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W413 N$825 N$826 "Straight Waveguide" sch_x=-3 sch_y=-10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W414 N$827 N$828 "Straight Waveguide" sch_x=-4 sch_y=-11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W415 N$829 N$830 "Straight Waveguide" sch_x=0 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W416 N$831 N$832 "Straight Waveguide" sch_x=-1 sch_y=-8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W417 N$833 N$834 "Straight Waveguide" sch_x=-1 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W418 N$835 N$836 "Straight Waveguide" sch_x=1 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W419 N$837 N$838 "Straight Waveguide" sch_x=1 sch_y=-8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W420 N$839 N$840 "Straight Waveguide" sch_x=0 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W421 N$841 N$842 "Straight Waveguide" sch_x=0 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W422 N$843 N$844 "Straight Waveguide" sch_x=-1 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W423 N$845 N$846 "Straight Waveguide" sch_x=-1 sch_y=-11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W424 N$847 N$848 "Straight Waveguide" sch_x=1 sch_y=-11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W425 N$849 N$850 "Straight Waveguide" sch_x=1 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W426 N$851 N$852 "Straight Waveguide" sch_x=0 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W427 N$853 N$854 "Straight Waveguide" sch_x=4 sch_y=-8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W428 N$855 N$856 "Straight Waveguide" sch_x=3 sch_y=-9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W429 N$857 N$858 "Straight Waveguide" sch_x=3 sch_y=-10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W430 N$859 N$860 "Straight Waveguide" sch_x=5 sch_y=-10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W431 N$861 N$862 "Straight Waveguide" sch_x=5 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W432 N$863 N$864 "Straight Waveguide" sch_x=4 sch_y=-11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W433 N$865 N$866 "Straight Waveguide" sch_x=-4 sch_y=-12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W434 N$867 N$868 "Straight Waveguide" sch_x=-5 sch_y=-13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W435 N$869 N$870 "Straight Waveguide" sch_x=-5 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W436 N$871 N$872 "Straight Waveguide" sch_x=-3 sch_y=-13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W437 N$873 N$874 "Straight Waveguide" sch_x=-3 sch_y=-14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W438 N$875 N$876 "Straight Waveguide" sch_x=-4 sch_y=-15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W439 N$877 N$878 "Straight Waveguide" sch_x=0 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W440 N$879 N$880 "Straight Waveguide" sch_x=-1 sch_y=-12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W441 N$881 N$882 "Straight Waveguide" sch_x=-1 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W442 N$883 N$884 "Straight Waveguide" sch_x=1 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W443 N$885 N$886 "Straight Waveguide" sch_x=1 sch_y=-12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W444 N$887 N$888 "Straight Waveguide" sch_x=0 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W445 N$889 N$890 "Straight Waveguide" sch_x=0 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W446 N$891 N$892 "Straight Waveguide" sch_x=-1 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W447 N$893 N$894 "Straight Waveguide" sch_x=-1 sch_y=-15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W448 N$895 N$896 "Straight Waveguide" sch_x=1 sch_y=-15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W449 N$897 N$898 "Straight Waveguide" sch_x=1 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W450 N$899 N$900 "Straight Waveguide" sch_x=0 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W451 N$901 N$902 "Straight Waveguide" sch_x=4 sch_y=-12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W452 N$903 N$904 "Straight Waveguide" sch_x=3 sch_y=-13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W453 N$905 N$906 "Straight Waveguide" sch_x=3 sch_y=-14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W454 N$907 N$908 "Straight Waveguide" sch_x=5 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W455 N$909 N$910 "Straight Waveguide" sch_x=5 sch_y=-13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W456 N$911 N$912 "Straight Waveguide" sch_x=4 sch_y=-15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W457 N$914 N$913 "Straight Waveguide" sch_x=-13 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W458 N$916 N$915 "Straight Waveguide" sch_x=-13 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W459 N$918 N$917 "Straight Waveguide" sch_x=-13 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W460 N$920 N$919 "Straight Waveguide" sch_x=-13 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W461 N$922 N$921 "Straight Waveguide" sch_x=-13 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W462 N$924 N$923 "Straight Waveguide" sch_x=-13 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W463 N$926 N$925 "Straight Waveguide" sch_x=-11 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W464 N$928 N$927 "Straight Waveguide" sch_x=-11 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W465 N$930 N$929 "Straight Waveguide" sch_x=-11 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W466 N$932 N$931 "Straight Waveguide" sch_x=-11 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W467 N$934 N$933 "Straight Waveguide" sch_x=-9 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W468 N$936 N$935 "Straight Waveguide" sch_x=-9 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W469 N$937 N$938 "Straight Waveguide" sch_x=-9 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W470 N$939 N$940 "Straight Waveguide" sch_x=-8 sch_y=-10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W471 N$941 N$942 "Straight Waveguide" sch_x=-7 sch_y=-11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W472 N$943 N$944 "Straight Waveguide" sch_x=-7 sch_y=-12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W473 N$945 N$946 "Straight Waveguide" sch_x=-8 sch_y=-13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W474 N$947 N$948 "Straight Waveguide" sch_x=-9 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W475 N$949 N$950 "Straight Waveguide" sch_x=-10 sch_y=-9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W476 N$951 N$952 "Straight Waveguide" sch_x=-10 sch_y=-14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W477 N$953 N$954 "Straight Waveguide" sch_x=13 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W478 N$955 N$956 "Straight Waveguide" sch_x=13 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W479 N$957 N$958 "Straight Waveguide" sch_x=13 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W480 N$959 N$960 "Straight Waveguide" sch_x=13 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W481 N$961 N$962 "Straight Waveguide" sch_x=13 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W482 N$963 N$964 "Straight Waveguide" sch_x=13 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W483 N$965 N$966 "Straight Waveguide" sch_x=11 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W484 N$967 N$968 "Straight Waveguide" sch_x=11 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W485 N$969 N$970 "Straight Waveguide" sch_x=11 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W486 N$971 N$972 "Straight Waveguide" sch_x=11 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W487 N$973 N$974 "Straight Waveguide" sch_x=9 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W488 N$975 N$976 "Straight Waveguide" sch_x=9 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W489 N$978 N$977 "Straight Waveguide" sch_x=9 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W490 N$980 N$979 "Straight Waveguide" sch_x=8 sch_y=-10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W491 N$982 N$981 "Straight Waveguide" sch_x=7 sch_y=-11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W492 N$984 N$983 "Straight Waveguide" sch_x=7 sch_y=-12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W493 N$986 N$985 "Straight Waveguide" sch_x=8 sch_y=-13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W494 N$988 N$987 "Straight Waveguide" sch_x=9 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W495 N$990 N$989 "Straight Waveguide" sch_x=10 sch_y=-9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W496 N$992 N$991 "Straight Waveguide" sch_x=10 sch_y=-14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W497 N$994 N$993 "Straight Waveguide" sch_x=-29 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W498 N$996 N$995 "Straight Waveguide" sch_x=-29 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W499 N$998 N$997 "Straight Waveguide" sch_x=-29 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W500 N$1000 N$999 "Straight Waveguide" sch_x=-29 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W501 N$1002 N$1001 "Straight Waveguide" sch_x=-29 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W502 N$1004 N$1003 "Straight Waveguide" sch_x=-29 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W503 N$1006 N$1005 "Straight Waveguide" sch_x=-29 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W504 N$1008 N$1007 "Straight Waveguide" sch_x=-29 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W505 N$1010 N$1009 "Straight Waveguide" sch_x=-29 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W506 N$1012 N$1011 "Straight Waveguide" sch_x=-29 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W507 N$1014 N$1013 "Straight Waveguide" sch_x=-29 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W508 N$1016 N$1015 "Straight Waveguide" sch_x=-29 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W509 N$1018 N$1017 "Straight Waveguide" sch_x=-29 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W510 N$1020 N$1019 "Straight Waveguide" sch_x=-29 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W511 N$1022 N$1021 "Straight Waveguide" sch_x=-27 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W512 N$1024 N$1023 "Straight Waveguide" sch_x=-27 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W513 N$1026 N$1025 "Straight Waveguide" sch_x=-27 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W514 N$1028 N$1027 "Straight Waveguide" sch_x=-27 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W515 N$1030 N$1029 "Straight Waveguide" sch_x=-27 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W516 N$1032 N$1031 "Straight Waveguide" sch_x=-27 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W517 N$1034 N$1033 "Straight Waveguide" sch_x=-27 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W518 N$1036 N$1035 "Straight Waveguide" sch_x=-27 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W519 N$1038 N$1037 "Straight Waveguide" sch_x=-27 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W520 N$1040 N$1039 "Straight Waveguide" sch_x=-27 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W521 N$1042 N$1041 "Straight Waveguide" sch_x=-27 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W522 N$1044 N$1043 "Straight Waveguide" sch_x=-27 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W523 N$1046 N$1045 "Straight Waveguide" sch_x=-25 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W524 N$1048 N$1047 "Straight Waveguide" sch_x=-25 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W525 N$1050 N$1049 "Straight Waveguide" sch_x=-25 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W526 N$1052 N$1051 "Straight Waveguide" sch_x=-25 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W527 N$1054 N$1053 "Straight Waveguide" sch_x=-25 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W528 N$1056 N$1055 "Straight Waveguide" sch_x=-25 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W529 N$1058 N$1057 "Straight Waveguide" sch_x=-25 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W530 N$1060 N$1059 "Straight Waveguide" sch_x=-25 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W531 N$1062 N$1061 "Straight Waveguide" sch_x=-25 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W532 N$1064 N$1063 "Straight Waveguide" sch_x=-25 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W533 N$1066 N$1065 "Straight Waveguide" sch_x=-23 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W534 N$1068 N$1067 "Straight Waveguide" sch_x=-23 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W535 N$1070 N$1069 "Straight Waveguide" sch_x=-23 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W536 N$1072 N$1071 "Straight Waveguide" sch_x=-23 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W537 N$1074 N$1073 "Straight Waveguide" sch_x=-23 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W538 N$1076 N$1075 "Straight Waveguide" sch_x=-23 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W539 N$1078 N$1077 "Straight Waveguide" sch_x=-23 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W540 N$1080 N$1079 "Straight Waveguide" sch_x=-23 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W541 N$1082 N$1081 "Straight Waveguide" sch_x=-21 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W542 N$1084 N$1083 "Straight Waveguide" sch_x=-21 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W543 N$1086 N$1085 "Straight Waveguide" sch_x=-21 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W544 N$1088 N$1087 "Straight Waveguide" sch_x=-21 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W545 N$1090 N$1089 "Straight Waveguide" sch_x=-21 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W546 N$1092 N$1091 "Straight Waveguide" sch_x=-21 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W547 N$1094 N$1093 "Straight Waveguide" sch_x=-19 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W548 N$1096 N$1095 "Straight Waveguide" sch_x=-19 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W549 N$1098 N$1097 "Straight Waveguide" sch_x=-19 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W550 N$1100 N$1099 "Straight Waveguide" sch_x=-19 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W551 N$1102 N$1101 "Straight Waveguide" sch_x=-17 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W552 N$1104 N$1103 "Straight Waveguide" sch_x=-17 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W553 N$1105 N$1106 "Straight Waveguide" sch_x=-21 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W554 N$1107 N$1108 "Straight Waveguide" sch_x=-20 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W555 N$1109 N$1110 "Straight Waveguide" sch_x=-19 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W556 N$1111 N$1112 "Straight Waveguide" sch_x=-18 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W557 N$1113 N$1114 "Straight Waveguide" sch_x=-17 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W558 N$1115 N$1116 "Straight Waveguide" sch_x=-16 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W559 N$1117 N$1118 "Straight Waveguide" sch_x=-15 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W560 N$1119 N$1120 "Straight Waveguide" sch_x=-15 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W561 N$1121 N$1122 "Straight Waveguide" sch_x=-16 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W562 N$1123 N$1124 "Straight Waveguide" sch_x=-17 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W563 N$1125 N$1126 "Straight Waveguide" sch_x=-18 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W564 N$1127 N$1128 "Straight Waveguide" sch_x=-19 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W565 N$1129 N$1130 "Straight Waveguide" sch_x=-20 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W566 N$1131 N$1132 "Straight Waveguide" sch_x=-21 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W567 N$1133 N$1134 "Straight Waveguide" sch_x=-22 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W568 N$1135 N$1136 "Straight Waveguide" sch_x=-22 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W569 N$1137 N$1138 "Straight Waveguide" sch_x=29 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W570 N$1139 N$1140 "Straight Waveguide" sch_x=29 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W571 N$1141 N$1142 "Straight Waveguide" sch_x=29 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W572 N$1143 N$1144 "Straight Waveguide" sch_x=29 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W573 N$1145 N$1146 "Straight Waveguide" sch_x=29 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W574 N$1147 N$1148 "Straight Waveguide" sch_x=29 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W575 N$1149 N$1150 "Straight Waveguide" sch_x=29 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W576 N$1151 N$1152 "Straight Waveguide" sch_x=29 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W577 N$1153 N$1154 "Straight Waveguide" sch_x=29 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W578 N$1155 N$1156 "Straight Waveguide" sch_x=29 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W579 N$1157 N$1158 "Straight Waveguide" sch_x=29 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W580 N$1159 N$1160 "Straight Waveguide" sch_x=29 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W581 N$1161 N$1162 "Straight Waveguide" sch_x=29 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W582 N$1163 N$1164 "Straight Waveguide" sch_x=29 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W583 N$1165 N$1166 "Straight Waveguide" sch_x=27 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W584 N$1167 N$1168 "Straight Waveguide" sch_x=27 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W585 N$1169 N$1170 "Straight Waveguide" sch_x=27 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W586 N$1171 N$1172 "Straight Waveguide" sch_x=27 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W587 N$1173 N$1174 "Straight Waveguide" sch_x=27 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W588 N$1175 N$1176 "Straight Waveguide" sch_x=27 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W589 N$1177 N$1178 "Straight Waveguide" sch_x=27 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W590 N$1179 N$1180 "Straight Waveguide" sch_x=27 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W591 N$1181 N$1182 "Straight Waveguide" sch_x=27 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W592 N$1183 N$1184 "Straight Waveguide" sch_x=27 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W593 N$1185 N$1186 "Straight Waveguide" sch_x=27 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W594 N$1187 N$1188 "Straight Waveguide" sch_x=27 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W595 N$1189 N$1190 "Straight Waveguide" sch_x=25 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W596 N$1191 N$1192 "Straight Waveguide" sch_x=25 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W597 N$1193 N$1194 "Straight Waveguide" sch_x=25 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W598 N$1195 N$1196 "Straight Waveguide" sch_x=25 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W599 N$1197 N$1198 "Straight Waveguide" sch_x=25 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W600 N$1199 N$1200 "Straight Waveguide" sch_x=25 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W601 N$1201 N$1202 "Straight Waveguide" sch_x=25 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W602 N$1203 N$1204 "Straight Waveguide" sch_x=25 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W603 N$1205 N$1206 "Straight Waveguide" sch_x=25 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W604 N$1207 N$1208 "Straight Waveguide" sch_x=25 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W605 N$1209 N$1210 "Straight Waveguide" sch_x=23 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W606 N$1211 N$1212 "Straight Waveguide" sch_x=23 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W607 N$1213 N$1214 "Straight Waveguide" sch_x=23 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W608 N$1215 N$1216 "Straight Waveguide" sch_x=23 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W609 N$1217 N$1218 "Straight Waveguide" sch_x=23 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W610 N$1219 N$1220 "Straight Waveguide" sch_x=23 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W611 N$1221 N$1222 "Straight Waveguide" sch_x=23 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W612 N$1223 N$1224 "Straight Waveguide" sch_x=23 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W613 N$1225 N$1226 "Straight Waveguide" sch_x=21 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W614 N$1227 N$1228 "Straight Waveguide" sch_x=21 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W615 N$1229 N$1230 "Straight Waveguide" sch_x=21 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W616 N$1231 N$1232 "Straight Waveguide" sch_x=21 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W617 N$1233 N$1234 "Straight Waveguide" sch_x=21 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W618 N$1235 N$1236 "Straight Waveguide" sch_x=21 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W619 N$1237 N$1238 "Straight Waveguide" sch_x=19 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W620 N$1239 N$1240 "Straight Waveguide" sch_x=19 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W621 N$1241 N$1242 "Straight Waveguide" sch_x=19 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W622 N$1243 N$1244 "Straight Waveguide" sch_x=19 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W623 N$1245 N$1246 "Straight Waveguide" sch_x=17 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W624 N$1247 N$1248 "Straight Waveguide" sch_x=17 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W625 N$1250 N$1249 "Straight Waveguide" sch_x=21 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W626 N$1252 N$1251 "Straight Waveguide" sch_x=20 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W627 N$1254 N$1253 "Straight Waveguide" sch_x=19 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W628 N$1256 N$1255 "Straight Waveguide" sch_x=18 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W629 N$1258 N$1257 "Straight Waveguide" sch_x=17 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W630 N$1260 N$1259 "Straight Waveguide" sch_x=16 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W631 N$1262 N$1261 "Straight Waveguide" sch_x=15 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W632 N$1264 N$1263 "Straight Waveguide" sch_x=15 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W633 N$1266 N$1265 "Straight Waveguide" sch_x=16 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W634 N$1268 N$1267 "Straight Waveguide" sch_x=17 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W635 N$1270 N$1269 "Straight Waveguide" sch_x=18 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W636 N$1272 N$1271 "Straight Waveguide" sch_x=19 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W637 N$1274 N$1273 "Straight Waveguide" sch_x=20 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W638 N$1276 N$1275 "Straight Waveguide" sch_x=21 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W639 N$1278 N$1277 "Straight Waveguide" sch_x=22 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W640 N$1280 N$1279 "Straight Waveguide" sch_x=22 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W641 N$1282 N$1281 "Straight Waveguide" sch_x=-61 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W642 N$1284 N$1283 "Straight Waveguide" sch_x=-61 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W643 N$1286 N$1285 "Straight Waveguide" sch_x=-61 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W644 N$1288 N$1287 "Straight Waveguide" sch_x=-61 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W645 N$1290 N$1289 "Straight Waveguide" sch_x=-61 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W646 N$1292 N$1291 "Straight Waveguide" sch_x=-61 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W647 N$1294 N$1293 "Straight Waveguide" sch_x=-61 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W648 N$1296 N$1295 "Straight Waveguide" sch_x=-61 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W649 N$1298 N$1297 "Straight Waveguide" sch_x=-61 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W650 N$1300 N$1299 "Straight Waveguide" sch_x=-61 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W651 N$1302 N$1301 "Straight Waveguide" sch_x=-61 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W652 N$1304 N$1303 "Straight Waveguide" sch_x=-61 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W653 N$1306 N$1305 "Straight Waveguide" sch_x=-61 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W654 N$1308 N$1307 "Straight Waveguide" sch_x=-61 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W655 N$1310 N$1309 "Straight Waveguide" sch_x=-61 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W656 N$1312 N$1311 "Straight Waveguide" sch_x=-61 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W657 N$1314 N$1313 "Straight Waveguide" sch_x=-61 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W658 N$1316 N$1315 "Straight Waveguide" sch_x=-61 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W659 N$1318 N$1317 "Straight Waveguide" sch_x=-61 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W660 N$1320 N$1319 "Straight Waveguide" sch_x=-61 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W661 N$1322 N$1321 "Straight Waveguide" sch_x=-61 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W662 N$1324 N$1323 "Straight Waveguide" sch_x=-61 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W663 N$1326 N$1325 "Straight Waveguide" sch_x=-61 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W664 N$1328 N$1327 "Straight Waveguide" sch_x=-61 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W665 N$1330 N$1329 "Straight Waveguide" sch_x=-61 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W666 N$1332 N$1331 "Straight Waveguide" sch_x=-61 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W667 N$1334 N$1333 "Straight Waveguide" sch_x=-61 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W668 N$1336 N$1335 "Straight Waveguide" sch_x=-61 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W669 N$1338 N$1337 "Straight Waveguide" sch_x=-61 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W670 N$1340 N$1339 "Straight Waveguide" sch_x=-61 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W671 N$1342 N$1341 "Straight Waveguide" sch_x=-59 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W672 N$1344 N$1343 "Straight Waveguide" sch_x=-59 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W673 N$1346 N$1345 "Straight Waveguide" sch_x=-59 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W674 N$1348 N$1347 "Straight Waveguide" sch_x=-59 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W675 N$1350 N$1349 "Straight Waveguide" sch_x=-59 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W676 N$1352 N$1351 "Straight Waveguide" sch_x=-59 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W677 N$1354 N$1353 "Straight Waveguide" sch_x=-59 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W678 N$1356 N$1355 "Straight Waveguide" sch_x=-59 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W679 N$1358 N$1357 "Straight Waveguide" sch_x=-59 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W680 N$1360 N$1359 "Straight Waveguide" sch_x=-59 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W681 N$1362 N$1361 "Straight Waveguide" sch_x=-59 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W682 N$1364 N$1363 "Straight Waveguide" sch_x=-59 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W683 N$1366 N$1365 "Straight Waveguide" sch_x=-59 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W684 N$1368 N$1367 "Straight Waveguide" sch_x=-59 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W685 N$1370 N$1369 "Straight Waveguide" sch_x=-59 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W686 N$1372 N$1371 "Straight Waveguide" sch_x=-59 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W687 N$1374 N$1373 "Straight Waveguide" sch_x=-59 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W688 N$1376 N$1375 "Straight Waveguide" sch_x=-59 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W689 N$1378 N$1377 "Straight Waveguide" sch_x=-59 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W690 N$1380 N$1379 "Straight Waveguide" sch_x=-59 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W691 N$1382 N$1381 "Straight Waveguide" sch_x=-59 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W692 N$1384 N$1383 "Straight Waveguide" sch_x=-59 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W693 N$1386 N$1385 "Straight Waveguide" sch_x=-59 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W694 N$1388 N$1387 "Straight Waveguide" sch_x=-59 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W695 N$1390 N$1389 "Straight Waveguide" sch_x=-59 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W696 N$1392 N$1391 "Straight Waveguide" sch_x=-59 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W697 N$1394 N$1393 "Straight Waveguide" sch_x=-59 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W698 N$1396 N$1395 "Straight Waveguide" sch_x=-59 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W699 N$1398 N$1397 "Straight Waveguide" sch_x=-57 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W700 N$1400 N$1399 "Straight Waveguide" sch_x=-57 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W701 N$1402 N$1401 "Straight Waveguide" sch_x=-57 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W702 N$1404 N$1403 "Straight Waveguide" sch_x=-57 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W703 N$1406 N$1405 "Straight Waveguide" sch_x=-57 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W704 N$1408 N$1407 "Straight Waveguide" sch_x=-57 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W705 N$1410 N$1409 "Straight Waveguide" sch_x=-57 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W706 N$1412 N$1411 "Straight Waveguide" sch_x=-57 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W707 N$1414 N$1413 "Straight Waveguide" sch_x=-57 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W708 N$1416 N$1415 "Straight Waveguide" sch_x=-57 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W709 N$1418 N$1417 "Straight Waveguide" sch_x=-57 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W710 N$1420 N$1419 "Straight Waveguide" sch_x=-57 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W711 N$1422 N$1421 "Straight Waveguide" sch_x=-57 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W712 N$1424 N$1423 "Straight Waveguide" sch_x=-57 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W713 N$1426 N$1425 "Straight Waveguide" sch_x=-57 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W714 N$1428 N$1427 "Straight Waveguide" sch_x=-57 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W715 N$1430 N$1429 "Straight Waveguide" sch_x=-57 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W716 N$1432 N$1431 "Straight Waveguide" sch_x=-57 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W717 N$1434 N$1433 "Straight Waveguide" sch_x=-57 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W718 N$1436 N$1435 "Straight Waveguide" sch_x=-57 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W719 N$1438 N$1437 "Straight Waveguide" sch_x=-57 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W720 N$1440 N$1439 "Straight Waveguide" sch_x=-57 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W721 N$1442 N$1441 "Straight Waveguide" sch_x=-57 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W722 N$1444 N$1443 "Straight Waveguide" sch_x=-57 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W723 N$1446 N$1445 "Straight Waveguide" sch_x=-57 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W724 N$1448 N$1447 "Straight Waveguide" sch_x=-57 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W725 N$1450 N$1449 "Straight Waveguide" sch_x=-55 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W726 N$1452 N$1451 "Straight Waveguide" sch_x=-55 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W727 N$1454 N$1453 "Straight Waveguide" sch_x=-55 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W728 N$1456 N$1455 "Straight Waveguide" sch_x=-55 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W729 N$1458 N$1457 "Straight Waveguide" sch_x=-55 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W730 N$1460 N$1459 "Straight Waveguide" sch_x=-55 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W731 N$1462 N$1461 "Straight Waveguide" sch_x=-55 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W732 N$1464 N$1463 "Straight Waveguide" sch_x=-55 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W733 N$1466 N$1465 "Straight Waveguide" sch_x=-55 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W734 N$1468 N$1467 "Straight Waveguide" sch_x=-55 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W735 N$1470 N$1469 "Straight Waveguide" sch_x=-55 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W736 N$1472 N$1471 "Straight Waveguide" sch_x=-55 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W737 N$1474 N$1473 "Straight Waveguide" sch_x=-55 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W738 N$1476 N$1475 "Straight Waveguide" sch_x=-55 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W739 N$1478 N$1477 "Straight Waveguide" sch_x=-55 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W740 N$1480 N$1479 "Straight Waveguide" sch_x=-55 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W741 N$1482 N$1481 "Straight Waveguide" sch_x=-55 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W742 N$1484 N$1483 "Straight Waveguide" sch_x=-55 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W743 N$1486 N$1485 "Straight Waveguide" sch_x=-55 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W744 N$1488 N$1487 "Straight Waveguide" sch_x=-55 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W745 N$1490 N$1489 "Straight Waveguide" sch_x=-55 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W746 N$1492 N$1491 "Straight Waveguide" sch_x=-55 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W747 N$1494 N$1493 "Straight Waveguide" sch_x=-55 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W748 N$1496 N$1495 "Straight Waveguide" sch_x=-55 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W749 N$1498 N$1497 "Straight Waveguide" sch_x=-53 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W750 N$1500 N$1499 "Straight Waveguide" sch_x=-53 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W751 N$1502 N$1501 "Straight Waveguide" sch_x=-53 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W752 N$1504 N$1503 "Straight Waveguide" sch_x=-53 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W753 N$1506 N$1505 "Straight Waveguide" sch_x=-53 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W754 N$1508 N$1507 "Straight Waveguide" sch_x=-53 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W755 N$1510 N$1509 "Straight Waveguide" sch_x=-53 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W756 N$1512 N$1511 "Straight Waveguide" sch_x=-53 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W757 N$1514 N$1513 "Straight Waveguide" sch_x=-53 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W758 N$1516 N$1515 "Straight Waveguide" sch_x=-53 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W759 N$1518 N$1517 "Straight Waveguide" sch_x=-53 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W760 N$1520 N$1519 "Straight Waveguide" sch_x=-53 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W761 N$1522 N$1521 "Straight Waveguide" sch_x=-53 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W762 N$1524 N$1523 "Straight Waveguide" sch_x=-53 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W763 N$1526 N$1525 "Straight Waveguide" sch_x=-53 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W764 N$1528 N$1527 "Straight Waveguide" sch_x=-53 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W765 N$1530 N$1529 "Straight Waveguide" sch_x=-53 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W766 N$1532 N$1531 "Straight Waveguide" sch_x=-53 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W767 N$1534 N$1533 "Straight Waveguide" sch_x=-53 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W768 N$1536 N$1535 "Straight Waveguide" sch_x=-53 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W769 N$1538 N$1537 "Straight Waveguide" sch_x=-53 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W770 N$1540 N$1539 "Straight Waveguide" sch_x=-53 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W771 N$1542 N$1541 "Straight Waveguide" sch_x=-51 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W772 N$1544 N$1543 "Straight Waveguide" sch_x=-51 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W773 N$1546 N$1545 "Straight Waveguide" sch_x=-51 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W774 N$1548 N$1547 "Straight Waveguide" sch_x=-51 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W775 N$1550 N$1549 "Straight Waveguide" sch_x=-51 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W776 N$1552 N$1551 "Straight Waveguide" sch_x=-51 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W777 N$1554 N$1553 "Straight Waveguide" sch_x=-51 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W778 N$1556 N$1555 "Straight Waveguide" sch_x=-51 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W779 N$1558 N$1557 "Straight Waveguide" sch_x=-51 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W780 N$1560 N$1559 "Straight Waveguide" sch_x=-51 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W781 N$1562 N$1561 "Straight Waveguide" sch_x=-51 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W782 N$1564 N$1563 "Straight Waveguide" sch_x=-51 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W783 N$1566 N$1565 "Straight Waveguide" sch_x=-51 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W784 N$1568 N$1567 "Straight Waveguide" sch_x=-51 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W785 N$1570 N$1569 "Straight Waveguide" sch_x=-51 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W786 N$1572 N$1571 "Straight Waveguide" sch_x=-51 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W787 N$1574 N$1573 "Straight Waveguide" sch_x=-51 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W788 N$1576 N$1575 "Straight Waveguide" sch_x=-51 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W789 N$1578 N$1577 "Straight Waveguide" sch_x=-51 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W790 N$1580 N$1579 "Straight Waveguide" sch_x=-51 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W791 N$1582 N$1581 "Straight Waveguide" sch_x=-49 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W792 N$1584 N$1583 "Straight Waveguide" sch_x=-49 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W793 N$1586 N$1585 "Straight Waveguide" sch_x=-49 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W794 N$1588 N$1587 "Straight Waveguide" sch_x=-49 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W795 N$1590 N$1589 "Straight Waveguide" sch_x=-49 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W796 N$1592 N$1591 "Straight Waveguide" sch_x=-49 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W797 N$1594 N$1593 "Straight Waveguide" sch_x=-49 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W798 N$1596 N$1595 "Straight Waveguide" sch_x=-49 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W799 N$1598 N$1597 "Straight Waveguide" sch_x=-49 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W800 N$1600 N$1599 "Straight Waveguide" sch_x=-49 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W801 N$1602 N$1601 "Straight Waveguide" sch_x=-49 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W802 N$1604 N$1603 "Straight Waveguide" sch_x=-49 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W803 N$1606 N$1605 "Straight Waveguide" sch_x=-49 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W804 N$1608 N$1607 "Straight Waveguide" sch_x=-49 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W805 N$1610 N$1609 "Straight Waveguide" sch_x=-49 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W806 N$1612 N$1611 "Straight Waveguide" sch_x=-49 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W807 N$1614 N$1613 "Straight Waveguide" sch_x=-49 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W808 N$1616 N$1615 "Straight Waveguide" sch_x=-49 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W809 N$1618 N$1617 "Straight Waveguide" sch_x=-47 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W810 N$1620 N$1619 "Straight Waveguide" sch_x=-47 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W811 N$1622 N$1621 "Straight Waveguide" sch_x=-47 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W812 N$1624 N$1623 "Straight Waveguide" sch_x=-47 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W813 N$1626 N$1625 "Straight Waveguide" sch_x=-47 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W814 N$1628 N$1627 "Straight Waveguide" sch_x=-47 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W815 N$1630 N$1629 "Straight Waveguide" sch_x=-47 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W816 N$1632 N$1631 "Straight Waveguide" sch_x=-47 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W817 N$1634 N$1633 "Straight Waveguide" sch_x=-47 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W818 N$1636 N$1635 "Straight Waveguide" sch_x=-47 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W819 N$1638 N$1637 "Straight Waveguide" sch_x=-47 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W820 N$1640 N$1639 "Straight Waveguide" sch_x=-47 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W821 N$1642 N$1641 "Straight Waveguide" sch_x=-47 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W822 N$1644 N$1643 "Straight Waveguide" sch_x=-47 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W823 N$1646 N$1645 "Straight Waveguide" sch_x=-47 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W824 N$1648 N$1647 "Straight Waveguide" sch_x=-47 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W825 N$1650 N$1649 "Straight Waveguide" sch_x=-45 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W826 N$1652 N$1651 "Straight Waveguide" sch_x=-45 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W827 N$1654 N$1653 "Straight Waveguide" sch_x=-45 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W828 N$1656 N$1655 "Straight Waveguide" sch_x=-45 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W829 N$1658 N$1657 "Straight Waveguide" sch_x=-45 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W830 N$1660 N$1659 "Straight Waveguide" sch_x=-45 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W831 N$1662 N$1661 "Straight Waveguide" sch_x=-45 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W832 N$1664 N$1663 "Straight Waveguide" sch_x=-45 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W833 N$1666 N$1665 "Straight Waveguide" sch_x=-45 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W834 N$1668 N$1667 "Straight Waveguide" sch_x=-45 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W835 N$1670 N$1669 "Straight Waveguide" sch_x=-45 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W836 N$1672 N$1671 "Straight Waveguide" sch_x=-45 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W837 N$1674 N$1673 "Straight Waveguide" sch_x=-45 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W838 N$1676 N$1675 "Straight Waveguide" sch_x=-45 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W839 N$1678 N$1677 "Straight Waveguide" sch_x=-43 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W840 N$1680 N$1679 "Straight Waveguide" sch_x=-43 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W841 N$1682 N$1681 "Straight Waveguide" sch_x=-43 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W842 N$1684 N$1683 "Straight Waveguide" sch_x=-43 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W843 N$1686 N$1685 "Straight Waveguide" sch_x=-43 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W844 N$1688 N$1687 "Straight Waveguide" sch_x=-43 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W845 N$1690 N$1689 "Straight Waveguide" sch_x=-43 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W846 N$1692 N$1691 "Straight Waveguide" sch_x=-43 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W847 N$1694 N$1693 "Straight Waveguide" sch_x=-43 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W848 N$1696 N$1695 "Straight Waveguide" sch_x=-43 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W849 N$1698 N$1697 "Straight Waveguide" sch_x=-43 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W850 N$1700 N$1699 "Straight Waveguide" sch_x=-43 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W851 N$1702 N$1701 "Straight Waveguide" sch_x=-41 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W852 N$1704 N$1703 "Straight Waveguide" sch_x=-41 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W853 N$1706 N$1705 "Straight Waveguide" sch_x=-41 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W854 N$1708 N$1707 "Straight Waveguide" sch_x=-41 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W855 N$1710 N$1709 "Straight Waveguide" sch_x=-41 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W856 N$1712 N$1711 "Straight Waveguide" sch_x=-41 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W857 N$1714 N$1713 "Straight Waveguide" sch_x=-41 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W858 N$1716 N$1715 "Straight Waveguide" sch_x=-41 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W859 N$1718 N$1717 "Straight Waveguide" sch_x=-41 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W860 N$1720 N$1719 "Straight Waveguide" sch_x=-41 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W861 N$1722 N$1721 "Straight Waveguide" sch_x=-39 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W862 N$1724 N$1723 "Straight Waveguide" sch_x=-39 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W863 N$1726 N$1725 "Straight Waveguide" sch_x=-39 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W864 N$1728 N$1727 "Straight Waveguide" sch_x=-39 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W865 N$1730 N$1729 "Straight Waveguide" sch_x=-39 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W866 N$1732 N$1731 "Straight Waveguide" sch_x=-39 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W867 N$1734 N$1733 "Straight Waveguide" sch_x=-39 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W868 N$1736 N$1735 "Straight Waveguide" sch_x=-39 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W869 N$1738 N$1737 "Straight Waveguide" sch_x=-37 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W870 N$1740 N$1739 "Straight Waveguide" sch_x=-37 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W871 N$1742 N$1741 "Straight Waveguide" sch_x=-37 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W872 N$1744 N$1743 "Straight Waveguide" sch_x=-37 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W873 N$1746 N$1745 "Straight Waveguide" sch_x=-37 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W874 N$1748 N$1747 "Straight Waveguide" sch_x=-37 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W875 N$1750 N$1749 "Straight Waveguide" sch_x=-35 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W876 N$1752 N$1751 "Straight Waveguide" sch_x=-35 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W877 N$1754 N$1753 "Straight Waveguide" sch_x=-35 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W878 N$1756 N$1755 "Straight Waveguide" sch_x=-35 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W879 N$1758 N$1757 "Straight Waveguide" sch_x=-33 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W880 N$1760 N$1759 "Straight Waveguide" sch_x=-33 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W881 N$1761 N$1762 "Straight Waveguide" sch_x=-45 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W882 N$1763 N$1764 "Straight Waveguide" sch_x=-44 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W883 N$1765 N$1766 "Straight Waveguide" sch_x=-43 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W884 N$1767 N$1768 "Straight Waveguide" sch_x=-42 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W885 N$1769 N$1770 "Straight Waveguide" sch_x=-41 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W886 N$1771 N$1772 "Straight Waveguide" sch_x=-40 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W887 N$1773 N$1774 "Straight Waveguide" sch_x=-39 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W888 N$1775 N$1776 "Straight Waveguide" sch_x=-38 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W889 N$1777 N$1778 "Straight Waveguide" sch_x=-37 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W890 N$1779 N$1780 "Straight Waveguide" sch_x=-36 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W891 N$1781 N$1782 "Straight Waveguide" sch_x=-35 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W892 N$1783 N$1784 "Straight Waveguide" sch_x=-34 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W893 N$1785 N$1786 "Straight Waveguide" sch_x=-33 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W894 N$1787 N$1788 "Straight Waveguide" sch_x=-32 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W895 N$1789 N$1790 "Straight Waveguide" sch_x=-31 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W896 N$1791 N$1792 "Straight Waveguide" sch_x=-31 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W897 N$1793 N$1794 "Straight Waveguide" sch_x=-32 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W898 N$1795 N$1796 "Straight Waveguide" sch_x=-33 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W899 N$1797 N$1798 "Straight Waveguide" sch_x=-34 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W900 N$1799 N$1800 "Straight Waveguide" sch_x=-35 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W901 N$1801 N$1802 "Straight Waveguide" sch_x=-36 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W902 N$1803 N$1804 "Straight Waveguide" sch_x=-37 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W903 N$1805 N$1806 "Straight Waveguide" sch_x=-38 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W904 N$1807 N$1808 "Straight Waveguide" sch_x=-39 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W905 N$1809 N$1810 "Straight Waveguide" sch_x=-40 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W906 N$1811 N$1812 "Straight Waveguide" sch_x=-41 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W907 N$1813 N$1814 "Straight Waveguide" sch_x=-42 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W908 N$1815 N$1816 "Straight Waveguide" sch_x=-43 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W909 N$1817 N$1818 "Straight Waveguide" sch_x=-44 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W910 N$1819 N$1820 "Straight Waveguide" sch_x=-45 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W911 N$1821 N$1822 "Straight Waveguide" sch_x=-46 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W912 N$1823 N$1824 "Straight Waveguide" sch_x=-46 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W913 N$1825 N$1826 "Straight Waveguide" sch_x=61 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W914 N$1827 N$1828 "Straight Waveguide" sch_x=61 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W915 N$1829 N$1830 "Straight Waveguide" sch_x=61 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W916 N$1831 N$1832 "Straight Waveguide" sch_x=61 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W917 N$1833 N$1834 "Straight Waveguide" sch_x=61 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W918 N$1835 N$1836 "Straight Waveguide" sch_x=61 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W919 N$1837 N$1838 "Straight Waveguide" sch_x=61 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W920 N$1839 N$1840 "Straight Waveguide" sch_x=61 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W921 N$1841 N$1842 "Straight Waveguide" sch_x=61 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W922 N$1843 N$1844 "Straight Waveguide" sch_x=61 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W923 N$1845 N$1846 "Straight Waveguide" sch_x=61 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W924 N$1847 N$1848 "Straight Waveguide" sch_x=61 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W925 N$1849 N$1850 "Straight Waveguide" sch_x=61 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W926 N$1851 N$1852 "Straight Waveguide" sch_x=61 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W927 N$1853 N$1854 "Straight Waveguide" sch_x=61 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W928 N$1855 N$1856 "Straight Waveguide" sch_x=61 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W929 N$1857 N$1858 "Straight Waveguide" sch_x=61 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W930 N$1859 N$1860 "Straight Waveguide" sch_x=61 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W931 N$1861 N$1862 "Straight Waveguide" sch_x=61 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W932 N$1863 N$1864 "Straight Waveguide" sch_x=61 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W933 N$1865 N$1866 "Straight Waveguide" sch_x=61 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W934 N$1867 N$1868 "Straight Waveguide" sch_x=61 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W935 N$1869 N$1870 "Straight Waveguide" sch_x=61 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W936 N$1871 N$1872 "Straight Waveguide" sch_x=61 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W937 N$1873 N$1874 "Straight Waveguide" sch_x=61 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W938 N$1875 N$1876 "Straight Waveguide" sch_x=61 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W939 N$1877 N$1878 "Straight Waveguide" sch_x=61 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W940 N$1879 N$1880 "Straight Waveguide" sch_x=61 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W941 N$1881 N$1882 "Straight Waveguide" sch_x=61 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W942 N$1883 N$1884 "Straight Waveguide" sch_x=61 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W943 N$1885 N$1886 "Straight Waveguide" sch_x=59 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W944 N$1887 N$1888 "Straight Waveguide" sch_x=59 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W945 N$1889 N$1890 "Straight Waveguide" sch_x=59 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W946 N$1891 N$1892 "Straight Waveguide" sch_x=59 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W947 N$1893 N$1894 "Straight Waveguide" sch_x=59 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W948 N$1895 N$1896 "Straight Waveguide" sch_x=59 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W949 N$1897 N$1898 "Straight Waveguide" sch_x=59 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W950 N$1899 N$1900 "Straight Waveguide" sch_x=59 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W951 N$1901 N$1902 "Straight Waveguide" sch_x=59 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W952 N$1903 N$1904 "Straight Waveguide" sch_x=59 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W953 N$1905 N$1906 "Straight Waveguide" sch_x=59 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W954 N$1907 N$1908 "Straight Waveguide" sch_x=59 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W955 N$1909 N$1910 "Straight Waveguide" sch_x=59 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W956 N$1911 N$1912 "Straight Waveguide" sch_x=59 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W957 N$1913 N$1914 "Straight Waveguide" sch_x=59 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W958 N$1915 N$1916 "Straight Waveguide" sch_x=59 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W959 N$1917 N$1918 "Straight Waveguide" sch_x=59 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W960 N$1919 N$1920 "Straight Waveguide" sch_x=59 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W961 N$1921 N$1922 "Straight Waveguide" sch_x=59 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W962 N$1923 N$1924 "Straight Waveguide" sch_x=59 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W963 N$1925 N$1926 "Straight Waveguide" sch_x=59 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W964 N$1927 N$1928 "Straight Waveguide" sch_x=59 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W965 N$1929 N$1930 "Straight Waveguide" sch_x=59 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W966 N$1931 N$1932 "Straight Waveguide" sch_x=59 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W967 N$1933 N$1934 "Straight Waveguide" sch_x=59 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W968 N$1935 N$1936 "Straight Waveguide" sch_x=59 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W969 N$1937 N$1938 "Straight Waveguide" sch_x=59 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W970 N$1939 N$1940 "Straight Waveguide" sch_x=59 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W971 N$1941 N$1942 "Straight Waveguide" sch_x=57 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W972 N$1943 N$1944 "Straight Waveguide" sch_x=57 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W973 N$1945 N$1946 "Straight Waveguide" sch_x=57 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W974 N$1947 N$1948 "Straight Waveguide" sch_x=57 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W975 N$1949 N$1950 "Straight Waveguide" sch_x=57 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W976 N$1951 N$1952 "Straight Waveguide" sch_x=57 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W977 N$1953 N$1954 "Straight Waveguide" sch_x=57 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W978 N$1955 N$1956 "Straight Waveguide" sch_x=57 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W979 N$1957 N$1958 "Straight Waveguide" sch_x=57 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W980 N$1959 N$1960 "Straight Waveguide" sch_x=57 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W981 N$1961 N$1962 "Straight Waveguide" sch_x=57 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W982 N$1963 N$1964 "Straight Waveguide" sch_x=57 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W983 N$1965 N$1966 "Straight Waveguide" sch_x=57 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W984 N$1967 N$1968 "Straight Waveguide" sch_x=57 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W985 N$1969 N$1970 "Straight Waveguide" sch_x=57 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W986 N$1971 N$1972 "Straight Waveguide" sch_x=57 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W987 N$1973 N$1974 "Straight Waveguide" sch_x=57 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W988 N$1975 N$1976 "Straight Waveguide" sch_x=57 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W989 N$1977 N$1978 "Straight Waveguide" sch_x=57 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W990 N$1979 N$1980 "Straight Waveguide" sch_x=57 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W991 N$1981 N$1982 "Straight Waveguide" sch_x=57 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W992 N$1983 N$1984 "Straight Waveguide" sch_x=57 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W993 N$1985 N$1986 "Straight Waveguide" sch_x=57 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W994 N$1987 N$1988 "Straight Waveguide" sch_x=57 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W995 N$1989 N$1990 "Straight Waveguide" sch_x=57 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W996 N$1991 N$1992 "Straight Waveguide" sch_x=57 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W997 N$1993 N$1994 "Straight Waveguide" sch_x=55 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W998 N$1995 N$1996 "Straight Waveguide" sch_x=55 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W999 N$1997 N$1998 "Straight Waveguide" sch_x=55 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1000 N$1999 N$2000 "Straight Waveguide" sch_x=55 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1001 N$2001 N$2002 "Straight Waveguide" sch_x=55 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1002 N$2003 N$2004 "Straight Waveguide" sch_x=55 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1003 N$2005 N$2006 "Straight Waveguide" sch_x=55 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1004 N$2007 N$2008 "Straight Waveguide" sch_x=55 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1005 N$2009 N$2010 "Straight Waveguide" sch_x=55 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1006 N$2011 N$2012 "Straight Waveguide" sch_x=55 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1007 N$2013 N$2014 "Straight Waveguide" sch_x=55 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1008 N$2015 N$2016 "Straight Waveguide" sch_x=55 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1009 N$2017 N$2018 "Straight Waveguide" sch_x=55 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1010 N$2019 N$2020 "Straight Waveguide" sch_x=55 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1011 N$2021 N$2022 "Straight Waveguide" sch_x=55 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1012 N$2023 N$2024 "Straight Waveguide" sch_x=55 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1013 N$2025 N$2026 "Straight Waveguide" sch_x=55 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1014 N$2027 N$2028 "Straight Waveguide" sch_x=55 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1015 N$2029 N$2030 "Straight Waveguide" sch_x=55 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1016 N$2031 N$2032 "Straight Waveguide" sch_x=55 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1017 N$2033 N$2034 "Straight Waveguide" sch_x=55 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1018 N$2035 N$2036 "Straight Waveguide" sch_x=55 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1019 N$2037 N$2038 "Straight Waveguide" sch_x=55 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1020 N$2039 N$2040 "Straight Waveguide" sch_x=55 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1021 N$2041 N$2042 "Straight Waveguide" sch_x=53 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1022 N$2043 N$2044 "Straight Waveguide" sch_x=53 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1023 N$2045 N$2046 "Straight Waveguide" sch_x=53 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1024 N$2047 N$2048 "Straight Waveguide" sch_x=53 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1025 N$2049 N$2050 "Straight Waveguide" sch_x=53 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1026 N$2051 N$2052 "Straight Waveguide" sch_x=53 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1027 N$2053 N$2054 "Straight Waveguide" sch_x=53 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1028 N$2055 N$2056 "Straight Waveguide" sch_x=53 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1029 N$2057 N$2058 "Straight Waveguide" sch_x=53 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1030 N$2059 N$2060 "Straight Waveguide" sch_x=53 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1031 N$2061 N$2062 "Straight Waveguide" sch_x=53 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1032 N$2063 N$2064 "Straight Waveguide" sch_x=53 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1033 N$2065 N$2066 "Straight Waveguide" sch_x=53 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1034 N$2067 N$2068 "Straight Waveguide" sch_x=53 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1035 N$2069 N$2070 "Straight Waveguide" sch_x=53 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1036 N$2071 N$2072 "Straight Waveguide" sch_x=53 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1037 N$2073 N$2074 "Straight Waveguide" sch_x=53 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1038 N$2075 N$2076 "Straight Waveguide" sch_x=53 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1039 N$2077 N$2078 "Straight Waveguide" sch_x=53 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1040 N$2079 N$2080 "Straight Waveguide" sch_x=53 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1041 N$2081 N$2082 "Straight Waveguide" sch_x=53 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1042 N$2083 N$2084 "Straight Waveguide" sch_x=53 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1043 N$2085 N$2086 "Straight Waveguide" sch_x=51 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1044 N$2087 N$2088 "Straight Waveguide" sch_x=51 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1045 N$2089 N$2090 "Straight Waveguide" sch_x=51 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1046 N$2091 N$2092 "Straight Waveguide" sch_x=51 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1047 N$2093 N$2094 "Straight Waveguide" sch_x=51 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1048 N$2095 N$2096 "Straight Waveguide" sch_x=51 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1049 N$2097 N$2098 "Straight Waveguide" sch_x=51 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1050 N$2099 N$2100 "Straight Waveguide" sch_x=51 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1051 N$2101 N$2102 "Straight Waveguide" sch_x=51 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1052 N$2103 N$2104 "Straight Waveguide" sch_x=51 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1053 N$2105 N$2106 "Straight Waveguide" sch_x=51 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1054 N$2107 N$2108 "Straight Waveguide" sch_x=51 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1055 N$2109 N$2110 "Straight Waveguide" sch_x=51 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1056 N$2111 N$2112 "Straight Waveguide" sch_x=51 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1057 N$2113 N$2114 "Straight Waveguide" sch_x=51 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1058 N$2115 N$2116 "Straight Waveguide" sch_x=51 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1059 N$2117 N$2118 "Straight Waveguide" sch_x=51 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1060 N$2119 N$2120 "Straight Waveguide" sch_x=51 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1061 N$2121 N$2122 "Straight Waveguide" sch_x=51 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1062 N$2123 N$2124 "Straight Waveguide" sch_x=51 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1063 N$2125 N$2126 "Straight Waveguide" sch_x=49 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1064 N$2127 N$2128 "Straight Waveguide" sch_x=49 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1065 N$2129 N$2130 "Straight Waveguide" sch_x=49 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1066 N$2131 N$2132 "Straight Waveguide" sch_x=49 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1067 N$2133 N$2134 "Straight Waveguide" sch_x=49 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1068 N$2135 N$2136 "Straight Waveguide" sch_x=49 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1069 N$2137 N$2138 "Straight Waveguide" sch_x=49 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1070 N$2139 N$2140 "Straight Waveguide" sch_x=49 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1071 N$2141 N$2142 "Straight Waveguide" sch_x=49 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1072 N$2143 N$2144 "Straight Waveguide" sch_x=49 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1073 N$2145 N$2146 "Straight Waveguide" sch_x=49 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1074 N$2147 N$2148 "Straight Waveguide" sch_x=49 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1075 N$2149 N$2150 "Straight Waveguide" sch_x=49 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1076 N$2151 N$2152 "Straight Waveguide" sch_x=49 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1077 N$2153 N$2154 "Straight Waveguide" sch_x=49 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1078 N$2155 N$2156 "Straight Waveguide" sch_x=49 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1079 N$2157 N$2158 "Straight Waveguide" sch_x=49 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1080 N$2159 N$2160 "Straight Waveguide" sch_x=49 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1081 N$2161 N$2162 "Straight Waveguide" sch_x=47 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1082 N$2163 N$2164 "Straight Waveguide" sch_x=47 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1083 N$2165 N$2166 "Straight Waveguide" sch_x=47 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1084 N$2167 N$2168 "Straight Waveguide" sch_x=47 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1085 N$2169 N$2170 "Straight Waveguide" sch_x=47 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1086 N$2171 N$2172 "Straight Waveguide" sch_x=47 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1087 N$2173 N$2174 "Straight Waveguide" sch_x=47 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1088 N$2175 N$2176 "Straight Waveguide" sch_x=47 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1089 N$2177 N$2178 "Straight Waveguide" sch_x=47 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1090 N$2179 N$2180 "Straight Waveguide" sch_x=47 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1091 N$2181 N$2182 "Straight Waveguide" sch_x=47 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1092 N$2183 N$2184 "Straight Waveguide" sch_x=47 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1093 N$2185 N$2186 "Straight Waveguide" sch_x=47 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1094 N$2187 N$2188 "Straight Waveguide" sch_x=47 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1095 N$2189 N$2190 "Straight Waveguide" sch_x=47 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1096 N$2191 N$2192 "Straight Waveguide" sch_x=47 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1097 N$2193 N$2194 "Straight Waveguide" sch_x=45 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1098 N$2195 N$2196 "Straight Waveguide" sch_x=45 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1099 N$2197 N$2198 "Straight Waveguide" sch_x=45 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1100 N$2199 N$2200 "Straight Waveguide" sch_x=45 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1101 N$2201 N$2202 "Straight Waveguide" sch_x=45 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1102 N$2203 N$2204 "Straight Waveguide" sch_x=45 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1103 N$2205 N$2206 "Straight Waveguide" sch_x=45 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1104 N$2207 N$2208 "Straight Waveguide" sch_x=45 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1105 N$2209 N$2210 "Straight Waveguide" sch_x=45 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1106 N$2211 N$2212 "Straight Waveguide" sch_x=45 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1107 N$2213 N$2214 "Straight Waveguide" sch_x=45 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1108 N$2215 N$2216 "Straight Waveguide" sch_x=45 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1109 N$2217 N$2218 "Straight Waveguide" sch_x=45 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1110 N$2219 N$2220 "Straight Waveguide" sch_x=45 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1111 N$2221 N$2222 "Straight Waveguide" sch_x=43 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1112 N$2223 N$2224 "Straight Waveguide" sch_x=43 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1113 N$2225 N$2226 "Straight Waveguide" sch_x=43 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1114 N$2227 N$2228 "Straight Waveguide" sch_x=43 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1115 N$2229 N$2230 "Straight Waveguide" sch_x=43 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1116 N$2231 N$2232 "Straight Waveguide" sch_x=43 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1117 N$2233 N$2234 "Straight Waveguide" sch_x=43 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1118 N$2235 N$2236 "Straight Waveguide" sch_x=43 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1119 N$2237 N$2238 "Straight Waveguide" sch_x=43 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1120 N$2239 N$2240 "Straight Waveguide" sch_x=43 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1121 N$2241 N$2242 "Straight Waveguide" sch_x=43 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1122 N$2243 N$2244 "Straight Waveguide" sch_x=43 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1123 N$2245 N$2246 "Straight Waveguide" sch_x=41 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1124 N$2247 N$2248 "Straight Waveguide" sch_x=41 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1125 N$2249 N$2250 "Straight Waveguide" sch_x=41 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1126 N$2251 N$2252 "Straight Waveguide" sch_x=41 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1127 N$2253 N$2254 "Straight Waveguide" sch_x=41 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1128 N$2255 N$2256 "Straight Waveguide" sch_x=41 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1129 N$2257 N$2258 "Straight Waveguide" sch_x=41 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1130 N$2259 N$2260 "Straight Waveguide" sch_x=41 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1131 N$2261 N$2262 "Straight Waveguide" sch_x=41 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1132 N$2263 N$2264 "Straight Waveguide" sch_x=41 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1133 N$2265 N$2266 "Straight Waveguide" sch_x=39 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1134 N$2267 N$2268 "Straight Waveguide" sch_x=39 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1135 N$2269 N$2270 "Straight Waveguide" sch_x=39 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1136 N$2271 N$2272 "Straight Waveguide" sch_x=39 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1137 N$2273 N$2274 "Straight Waveguide" sch_x=39 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1138 N$2275 N$2276 "Straight Waveguide" sch_x=39 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1139 N$2277 N$2278 "Straight Waveguide" sch_x=39 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1140 N$2279 N$2280 "Straight Waveguide" sch_x=39 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1141 N$2281 N$2282 "Straight Waveguide" sch_x=37 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1142 N$2283 N$2284 "Straight Waveguide" sch_x=37 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1143 N$2285 N$2286 "Straight Waveguide" sch_x=37 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1144 N$2287 N$2288 "Straight Waveguide" sch_x=37 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1145 N$2289 N$2290 "Straight Waveguide" sch_x=37 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1146 N$2291 N$2292 "Straight Waveguide" sch_x=37 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1147 N$2293 N$2294 "Straight Waveguide" sch_x=35 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1148 N$2295 N$2296 "Straight Waveguide" sch_x=35 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1149 N$2297 N$2298 "Straight Waveguide" sch_x=35 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1150 N$2299 N$2300 "Straight Waveguide" sch_x=35 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1151 N$2301 N$2302 "Straight Waveguide" sch_x=33 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1152 N$2303 N$2304 "Straight Waveguide" sch_x=33 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1153 N$2306 N$2305 "Straight Waveguide" sch_x=45 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1154 N$2308 N$2307 "Straight Waveguide" sch_x=44 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1155 N$2310 N$2309 "Straight Waveguide" sch_x=43 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1156 N$2312 N$2311 "Straight Waveguide" sch_x=42 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1157 N$2314 N$2313 "Straight Waveguide" sch_x=41 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1158 N$2316 N$2315 "Straight Waveguide" sch_x=40 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1159 N$2318 N$2317 "Straight Waveguide" sch_x=39 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1160 N$2320 N$2319 "Straight Waveguide" sch_x=38 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1161 N$2322 N$2321 "Straight Waveguide" sch_x=37 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1162 N$2324 N$2323 "Straight Waveguide" sch_x=36 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1163 N$2326 N$2325 "Straight Waveguide" sch_x=35 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1164 N$2328 N$2327 "Straight Waveguide" sch_x=34 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1165 N$2330 N$2329 "Straight Waveguide" sch_x=33 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1166 N$2332 N$2331 "Straight Waveguide" sch_x=32 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1167 N$2334 N$2333 "Straight Waveguide" sch_x=31 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1168 N$2336 N$2335 "Straight Waveguide" sch_x=31 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1169 N$2338 N$2337 "Straight Waveguide" sch_x=32 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1170 N$2340 N$2339 "Straight Waveguide" sch_x=33 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1171 N$2342 N$2341 "Straight Waveguide" sch_x=34 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1172 N$2344 N$2343 "Straight Waveguide" sch_x=35 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1173 N$2346 N$2345 "Straight Waveguide" sch_x=36 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1174 N$2348 N$2347 "Straight Waveguide" sch_x=37 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1175 N$2350 N$2349 "Straight Waveguide" sch_x=38 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1176 N$2352 N$2351 "Straight Waveguide" sch_x=39 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1177 N$2354 N$2353 "Straight Waveguide" sch_x=40 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1178 N$2356 N$2355 "Straight Waveguide" sch_x=41 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1179 N$2358 N$2357 "Straight Waveguide" sch_x=42 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1180 N$2360 N$2359 "Straight Waveguide" sch_x=43 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1181 N$2362 N$2361 "Straight Waveguide" sch_x=44 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1182 N$2364 N$2363 "Straight Waveguide" sch_x=45 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1183 N$2366 N$2365 "Straight Waveguide" sch_x=46 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1184 N$2368 N$2367 "Straight Waveguide" sch_x=46 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
.ends HDBE
* - ONA
.ona input_unit=wavelength input_parameter=center_and_range center=1550e-9
  + range=100e-9 number_of_points=100 
  + minimum_loss=200
  + sensitivity=-200 
  + analysis_type=scattering_data
  + multithreading=user_defined number_of_threads=1 
 + input(1)=HDBE,N$2465
+ input(2)=HDBE,N$2467
+ input(3)=HDBE,N$2469
+ input(4)=HDBE,N$2471
+ input(5)=HDBE,N$2473
+ input(6)=HDBE,N$2475
+ input(7)=HDBE,N$2477
+ input(8)=HDBE,N$2479
+ input(9)=HDBE,N$2481
+ input(10)=HDBE,N$2483
+ input(11)=HDBE,N$2485
+ input(12)=HDBE,N$2487
+ input(13)=HDBE,N$2489
+ input(14)=HDBE,N$2491
+ input(15)=HDBE,N$2493
+ input(16)=HDBE,N$2495
  + output=HDBE,N$2369

HDBE  N$2369 N$2371 N$2373 N$2375 N$2377 N$2379 N$2381 N$2383 N$2385 N$2387 N$2389 N$2391 N$2393 N$2395 N$2397 N$2399 N$2465 N$2467 N$2469 N$2471 N$2473 N$2475 N$2477 N$2479 N$2481 N$2483 N$2485 N$2487 N$2489 N$2491 N$2493 N$2495 HDBE sch_x=0 sch_y=0
*
.end